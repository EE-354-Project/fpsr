module gandhi_up_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin

		if(({row_reg, col_reg}>=12'b000000000000) && ({row_reg, col_reg}<12'b000001011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b000001011100)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b000001011101) && ({row_reg, col_reg}<12'b000010010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b000010010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b000010010001) && ({row_reg, col_reg}<12'b000010010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b000010010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b000010010110) && ({row_reg, col_reg}<12'b000010011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b000010011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b000010011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b000010011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b000010011011) && ({row_reg, col_reg}<12'b000010011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b000010011111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b000010100000) && ({row_reg, col_reg}<12'b000011010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b000011010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b000011010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000011010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b000011010101) && ({row_reg, col_reg}<12'b000011011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b000011011000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b000011011001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=12'b000011011010) && ({row_reg, col_reg}<12'b000011011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000011011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000011011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b000011011110) && ({row_reg, col_reg}<12'b000011100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b000011100000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b000011100001) && ({row_reg, col_reg}<12'b000100010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b000100010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b000100010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b000100010010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b000100010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b000100010100) && ({row_reg, col_reg}<12'b000100010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000100010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b000100010111) && ({row_reg, col_reg}<12'b000100011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000100011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b000100011011) && ({row_reg, col_reg}<12'b000100011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000100011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b000100011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b000100011111)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=12'b000100100000) && ({row_reg, col_reg}<12'b000101001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b000101001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000101010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b000101010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b000101010011) && ({row_reg, col_reg}<12'b000101010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000101010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b000101010110) && ({row_reg, col_reg}<12'b000101011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000101011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b000101011010) && ({row_reg, col_reg}<12'b000101011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000101011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b000101011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000101011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000101011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b000101100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000101100001)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=12'b000101100010) && ({row_reg, col_reg}<12'b000110001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b000110001110) && ({row_reg, col_reg}<12'b000110010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000110010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b000110010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000110010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000110010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b000110010101) && ({row_reg, col_reg}<12'b000110010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b000110010111) && ({row_reg, col_reg}<12'b000110011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000110011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b000110011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b000110011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b000110011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000110011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000110011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000110011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000110100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000110100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b000110100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b000110100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b000110100100)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b000110100101) && ({row_reg, col_reg}<12'b000111001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b000111001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000111001110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b000111001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b000111010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000111010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b000111010010) && ({row_reg, col_reg}<12'b000111010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000111010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b000111010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000111011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b000111011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b000111011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000111011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000111011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b000111011101) && ({row_reg, col_reg}<12'b000111011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b000111011111) && ({row_reg, col_reg}<12'b000111100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000111100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b000111100010)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b000111100011)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=12'b000111100100) && ({row_reg, col_reg}<12'b001000001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001000001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001000001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=12'b001000001110) && ({row_reg, col_reg}<12'b001000010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b001000010010) && ({row_reg, col_reg}<12'b001000010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001000010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b001000010101) && ({row_reg, col_reg}<12'b001000011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001000011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b001000011010) && ({row_reg, col_reg}<12'b001000011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001000011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b001000011101) && ({row_reg, col_reg}<12'b001000011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001000011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b001000100000) && ({row_reg, col_reg}<12'b001000100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001000100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001000100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001000100100)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=12'b001000100101) && ({row_reg, col_reg}<12'b001001001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001001001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b001001001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001001001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001001001100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==12'b001001001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b001001001110) && ({row_reg, col_reg}<12'b001001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001001010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001001010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001001010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001001011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001001011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001001011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001001011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001001011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b001001011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b001001011110) && ({row_reg, col_reg}<12'b001001100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001001100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001001100100)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b001001100101) && ({row_reg, col_reg}<12'b001010001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b001010001011) && ({row_reg, col_reg}<12'b001010001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001010001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b001010001110) && ({row_reg, col_reg}<12'b001010010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001010010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001010010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001010010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b001010010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b001010010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001010010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001010011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001010011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001010011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b001010011011) && ({row_reg, col_reg}<12'b001010100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001010100101)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=12'b001010100110) && ({row_reg, col_reg}<12'b001011001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001011001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b001011001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b001011001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b001011001101) && ({row_reg, col_reg}<12'b001011001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001011001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001011010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001011010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b001011010010) && ({row_reg, col_reg}<12'b001011010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001011010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001011010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b001011010111) && ({row_reg, col_reg}<12'b001011011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b001011011001) && ({row_reg, col_reg}<12'b001011100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001011100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b001011100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001011100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b001011100101)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b001011100110) && ({row_reg, col_reg}<12'b001100001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001100001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b001100001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b001100001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001100001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001100001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001100001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001100010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001100010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001100010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b001100010011) && ({row_reg, col_reg}<12'b001100010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001100010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b001100010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001100010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b001100011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001100011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b001100011010) && ({row_reg, col_reg}<12'b001100100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001100100110)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=12'b001100100111) && ({row_reg, col_reg}<12'b001101001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001101001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001101001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b001101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001101001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b001101010001) && ({row_reg, col_reg}<12'b001101010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001101010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001101010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001101010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b001101011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001101011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b001101011010) && ({row_reg, col_reg}<12'b001101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001101100101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b001101100110)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}>=12'b001101100111) && ({row_reg, col_reg}<12'b001110001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001110001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001110001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001110001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001110001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b001110001110) && ({row_reg, col_reg}<12'b001110010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001110010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b001110010010) && ({row_reg, col_reg}<12'b001110010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001110010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001110010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001110010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001110010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b001110011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001110011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b001110011010) && ({row_reg, col_reg}<12'b001110011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001110011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b001110011111) && ({row_reg, col_reg}<12'b001110100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b001110100001) && ({row_reg, col_reg}<12'b001110100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b001110100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b001110100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001110100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b001110100110)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=12'b001110100111) && ({row_reg, col_reg}<12'b001111001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001111001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001111001011)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==12'b001111001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001111001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001111001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b001111001111) && ({row_reg, col_reg}<12'b001111010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b001111010001) && ({row_reg, col_reg}<12'b001111010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b001111010011) && ({row_reg, col_reg}<12'b001111010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001111010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b001111010110) && ({row_reg, col_reg}<12'b001111011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001111011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001111011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b001111011010) && ({row_reg, col_reg}<12'b001111011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001111011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b001111011111) && ({row_reg, col_reg}<12'b001111100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001111100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001111100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001111100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001111100111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b001111101000) && ({row_reg, col_reg}<12'b010000001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010000001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010000001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=12'b010000001100) && ({row_reg, col_reg}<12'b010000001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010000001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010000001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b010000010000) && ({row_reg, col_reg}<12'b010000010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010000010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010000010011) && ({row_reg, col_reg}<12'b010000010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010000010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b010000010110) && ({row_reg, col_reg}<12'b010000011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010000011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010000011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b010000011010) && ({row_reg, col_reg}<12'b010000011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010000011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b010000011101) && ({row_reg, col_reg}<12'b010000100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b010000100010) && ({row_reg, col_reg}<12'b010000100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010000100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b010000100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010000100111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b010000101000) && ({row_reg, col_reg}<12'b010001001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010001001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b010001001011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010001001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b010001001101) && ({row_reg, col_reg}<12'b010001001111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b010001001111) && ({row_reg, col_reg}<12'b010001010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010001010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010001010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b010001010110) && ({row_reg, col_reg}<12'b010001011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010001011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010001011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b010001011010) && ({row_reg, col_reg}<12'b010001011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b010001011111) && ({row_reg, col_reg}<12'b010001100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b010001100001) && ({row_reg, col_reg}<12'b010001100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b010001100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b010001100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010001100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b010001100110)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=12'b010001100111) && ({row_reg, col_reg}<12'b010010001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010010001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010010001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010010001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b010010001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b010010001110) && ({row_reg, col_reg}<12'b010010010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010010010000) && ({row_reg, col_reg}<12'b010010010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010010010011)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010010010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010010010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b010010010110) && ({row_reg, col_reg}<12'b010010011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010010011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010010011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b010010011010) && ({row_reg, col_reg}<12'b010010100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010010100111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b010010101000) && ({row_reg, col_reg}<12'b010011001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010011001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b010011001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010011001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010011001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010011001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010011001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b010011001111) && ({row_reg, col_reg}<12'b010011010001)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010011010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b010011010010) && ({row_reg, col_reg}<12'b010011010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010011010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010011010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010011010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b010011010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010011011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010011011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b010011011010) && ({row_reg, col_reg}<12'b010011100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010011100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010011100111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b010011101000) && ({row_reg, col_reg}<12'b010100001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010100001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b010100001010) && ({row_reg, col_reg}<12'b010100001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010100001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010100001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010100001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010100001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b010100010000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b010100010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010100010010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010100010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b010100010100) && ({row_reg, col_reg}<12'b010100010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010100010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b010100011000) && ({row_reg, col_reg}<12'b010100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010100011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010100011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010100011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010100011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b010100011110) && ({row_reg, col_reg}<12'b010100100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010100100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b010100100010) && ({row_reg, col_reg}<12'b010100100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010100100111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=12'b010100101000) && ({row_reg, col_reg}<12'b010101001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010101001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b010101001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010101001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010101001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b010101010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010101010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010101010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010101010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010101010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010101010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b010101010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010101011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b010101011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010101011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010101011011) && ({row_reg, col_reg}<12'b010101011101)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}>=12'b010101011101) && ({row_reg, col_reg}<12'b010101011111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010101011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010101100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010101100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010101100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b010101100011) && ({row_reg, col_reg}<12'b010101100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b010101100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010101100110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010101100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b010101101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b010101101001) && ({row_reg, col_reg}<12'b010101101011)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b010101101011) && ({row_reg, col_reg}<12'b010110001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b010110001001) && ({row_reg, col_reg}<12'b010110001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010110001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010110001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010110001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b010110001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010110001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b010110010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010110010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010110010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010110010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b010110010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010110010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010110010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010110011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b010110011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b010110011010) && ({row_reg, col_reg}<12'b010110011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010110011100) && ({row_reg, col_reg}<12'b010110011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010110011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010110011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010110100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b010110100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010110100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b010110100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010110100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010110100101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010110100110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b010110100111)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=12'b010110101000) && ({row_reg, col_reg}<12'b010111001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010111001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b010111001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010111001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b010111001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010111001101) && ({row_reg, col_reg}<12'b010111001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010111001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b010111010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010111010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010111010011) && ({row_reg, col_reg}<12'b010111010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010111010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b010111010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010111011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b010111011010) && ({row_reg, col_reg}<12'b010111011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010111011100) && ({row_reg, col_reg}<12'b010111011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010111011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b010111011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010111100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010111100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b010111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010111100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b010111100101) && ({row_reg, col_reg}<12'b010111100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010111100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010111101000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010111101001)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=12'b010111101010) && ({row_reg, col_reg}<12'b011000001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011000001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011000001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011000001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011000001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011000010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b011000010001) && ({row_reg, col_reg}<12'b011000010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b011000010011) && ({row_reg, col_reg}<12'b011000010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011000010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011000010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011000011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b011000011001) && ({row_reg, col_reg}<12'b011000011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011000011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011000011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011000011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011000011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011000011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b011000100000) && ({row_reg, col_reg}<12'b011000100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011000100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b011000100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011000100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011000100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011000100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011000101001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011000101010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b011000101011) && ({row_reg, col_reg}<12'b011001001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b011001001010) && ({row_reg, col_reg}<12'b011001001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011001001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011001001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011001001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b011001010000) && ({row_reg, col_reg}<12'b011001010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011001010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011001010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b011001010100) && ({row_reg, col_reg}<12'b011001010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011001010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b011001010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011001011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011001011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b011001011011) && ({row_reg, col_reg}<12'b011001011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011001011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011001011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011001011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011001100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011001100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011001100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011001100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011001100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011001100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b011001100110) && ({row_reg, col_reg}<12'b011001101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011001101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011001101001)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=12'b011001101010) && ({row_reg, col_reg}<12'b011010001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011010001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011010001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011010001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011010001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011010001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011010001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b011010010000) && ({row_reg, col_reg}<12'b011010010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011010010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011010010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b011010010101) && ({row_reg, col_reg}<12'b011010010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011010010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011010011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011010011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011010011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b011010011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011010011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011010011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011010011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011010011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b011010100000) && ({row_reg, col_reg}<12'b011010100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011010100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011010100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011010100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011010100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011010100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011010100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011010101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b011010101001) && ({row_reg, col_reg}<12'b011010101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011010101111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b011010110000) && ({row_reg, col_reg}<12'b011011001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011011001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011011001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011011001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b011011001110) && ({row_reg, col_reg}<12'b011011010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011011010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b011011010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011011010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011011010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011011010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b011011010101) && ({row_reg, col_reg}<12'b011011011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011011011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011011011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011011011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b011011011011) && ({row_reg, col_reg}<12'b011011011101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b011011011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011011011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011011011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b011011100000) && ({row_reg, col_reg}<12'b011011100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011011100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b011011100011) && ({row_reg, col_reg}<12'b011011100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011011100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011011100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011011100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011011101000)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=12'b011011101001) && ({row_reg, col_reg}<12'b011100001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011100001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011100001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b011100001101) && ({row_reg, col_reg}<12'b011100001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b011100001111) && ({row_reg, col_reg}<12'b011100010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011100010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011100010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011100010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011100010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b011100010101) && ({row_reg, col_reg}<12'b011100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011100011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011100011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011100011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011100011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011100011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011100011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b011100011111) && ({row_reg, col_reg}<12'b011100100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011100100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011100100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b011100100100) && ({row_reg, col_reg}<12'b011100100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011100100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011100100111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=12'b011100101000) && ({row_reg, col_reg}<12'b011101001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011101001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b011101001010) && ({row_reg, col_reg}<12'b011101001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011101001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011101001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011101001111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011101010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b011101010001) && ({row_reg, col_reg}<12'b011101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011101010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011101010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011101010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b011101010110) && ({row_reg, col_reg}<12'b011101011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011101011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011101011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011101011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011101011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b011101100000) && ({row_reg, col_reg}<12'b011101100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011101100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011101100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b011101100100) && ({row_reg, col_reg}<12'b011101100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b011101100110) && ({row_reg, col_reg}<12'b011101101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011101101000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b011101101001) && ({row_reg, col_reg}<12'b011110001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011110001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b011110001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011110001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011110001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011110010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011110010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011110010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011110010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011110010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b011110010110) && ({row_reg, col_reg}<12'b011110011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011110011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011110011100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b011110011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011110011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b011110011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b011110100000) && ({row_reg, col_reg}<12'b011110100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011110100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011110100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011110100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011110100101)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=12'b011110100110) && ({row_reg, col_reg}<12'b011111001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011111001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011111001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011111001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011111001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011111010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b011111010001) && ({row_reg, col_reg}<12'b011111010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011111010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011111010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b011111010110) && ({row_reg, col_reg}<12'b011111011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011111011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011111011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011111011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011111011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b011111011101) && ({row_reg, col_reg}<12'b011111011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b011111011111) && ({row_reg, col_reg}<12'b011111100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011111100010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b011111100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011111100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b011111100101) && ({row_reg, col_reg}<12'b011111101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011111101110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b011111101111) && ({row_reg, col_reg}<12'b100000001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b100000001011) && ({row_reg, col_reg}<12'b100000001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100000001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100000001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100000001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100000010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100000010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100000010010) && ({row_reg, col_reg}<12'b100000010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100000010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100000010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b100000010110) && ({row_reg, col_reg}<12'b100000011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100000011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100000011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100000011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b100000011011) && ({row_reg, col_reg}<12'b100000011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100000011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100000011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100000011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100000100000) && ({row_reg, col_reg}<12'b100000100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100000100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100000100011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b100000100100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=12'b100000100101) && ({row_reg, col_reg}<12'b100001000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b100001000010) && ({row_reg, col_reg}<12'b100001000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b100001000101) && ({row_reg, col_reg}<12'b100001001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100001001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100001001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b100001001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100001001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100001010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100001010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100001010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100001010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100001010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100001011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100001011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b100001011010) && ({row_reg, col_reg}<12'b100001011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100001100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100001100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b100001100010) && ({row_reg, col_reg}<12'b100001100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100001100100) && ({row_reg, col_reg}<12'b100001100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001100110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b100001100111) && ({row_reg, col_reg}<12'b100010001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100010001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100010001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100010001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100010001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100010001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100010001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100010001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100010010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b100010010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100010010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100010010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b100010010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100010010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100010010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100010010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100010011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100010011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100010011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100010011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100010011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100010011101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b100010011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100010011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100010100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100010100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100010100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b100010100011)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b100010100100) && ({row_reg, col_reg}<12'b100011000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100011000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100011001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100011001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100011001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100011001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100011001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100011001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100011001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100011001111) && ({row_reg, col_reg}<12'b100011010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b100011010001) && ({row_reg, col_reg}<12'b100011010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100011010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100011010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b100011010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100011010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100011010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b100011011000) && ({row_reg, col_reg}<12'b100011011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100011011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100011011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100011011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b100011011101) && ({row_reg, col_reg}<12'b100011100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100011100000) && ({row_reg, col_reg}<12'b100011100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100011100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100011100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100011100100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=12'b100011100101) && ({row_reg, col_reg}<12'b100100000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100100000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100100001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100100001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100100001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100100001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b100100001100) && ({row_reg, col_reg}<12'b100100001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100100001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100100001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100100010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100100010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100100010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100100010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100100010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100100010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b100100010110) && ({row_reg, col_reg}<12'b100100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b100100011001) && ({row_reg, col_reg}<12'b100100011011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100100011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100100011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100100011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100100100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b100100100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100100100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100100100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b100100100100) && ({row_reg, col_reg}<12'b100100100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100100100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b100100100111) && ({row_reg, col_reg}<12'b100100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100100101011)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b100100101100) && ({row_reg, col_reg}<12'b100101000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100101000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b100101000010) && ({row_reg, col_reg}<12'b100101000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100101000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100101000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100101000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b100101000111) && ({row_reg, col_reg}<12'b100101001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100101001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b100101001100) && ({row_reg, col_reg}<12'b100101001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100101001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100101010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b100101010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100101010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100101010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100101010110) && ({row_reg, col_reg}<12'b100101011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100101011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100101011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100101011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100101011100) && ({row_reg, col_reg}<12'b100101011110)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=12'b100101011110) && ({row_reg, col_reg}<12'b100101100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100101100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100101100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b100101100010) && ({row_reg, col_reg}<12'b100101100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100101100101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100101100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100101100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100101101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100101101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b100101101010) && ({row_reg, col_reg}<12'b100101101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100101101110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b100101101111) && ({row_reg, col_reg}<12'b100110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100110000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100110000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100110000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b100110000110) && ({row_reg, col_reg}<12'b100110001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100110001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100110001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100110001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100110001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b100110001100) && ({row_reg, col_reg}<12'b100110001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100110001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100110010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100110010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100110010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100110010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100110010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100110010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100110010111) && ({row_reg, col_reg}<12'b100110011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b100110011001) && ({row_reg, col_reg}<12'b100110011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b100110011100) && ({row_reg, col_reg}<12'b100110011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b100110011110) && ({row_reg, col_reg}<12'b100110100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100110100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100110100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100110100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100110100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b100110100100) && ({row_reg, col_reg}<12'b100110100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100110100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100110101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100110101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100110101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100110101011)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=12'b100110101100) && ({row_reg, col_reg}<12'b100111000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100111000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100111000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100111001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100111001001) && ({row_reg, col_reg}<12'b100111001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100111001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100111001100) && ({row_reg, col_reg}<12'b100111010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100111010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b100111010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b100111010010) && ({row_reg, col_reg}<12'b100111010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100111010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b100111010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100111010110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b100111010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100111011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b100111011001) && ({row_reg, col_reg}<12'b100111011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100111011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100111011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b100111100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100111100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100111100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b100111100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100111100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100111100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100111100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b100111100111) && ({row_reg, col_reg}<12'b100111101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100111101010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b100111101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100111101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100111101101)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=12'b100111101110) && ({row_reg, col_reg}<12'b101000000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101000000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101000000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101000000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b101000001000) && ({row_reg, col_reg}<12'b101000001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101000001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101000001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b101000001101) && ({row_reg, col_reg}<12'b101000010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101000010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101000010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101000010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101000010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101000010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b101000010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101000010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101000011000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b101000011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101000011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101000011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101000011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b101000011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101000011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b101000011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101000100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101000100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b101000100010) && ({row_reg, col_reg}<12'b101000100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101000100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b101000100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101000100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101000101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b101000101010) && ({row_reg, col_reg}<12'b101000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101000101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101000101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101000101110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b101000101111) && ({row_reg, col_reg}<12'b101001000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101001000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101001000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101001000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101001000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101001001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101001001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101001001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101001001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101001001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b101001001101) && ({row_reg, col_reg}<12'b101001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101001010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101001010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b101001010011) && ({row_reg, col_reg}<12'b101001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101001010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101001010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101001011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b101001011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101001011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101001011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101001011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101001011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b101001011110) && ({row_reg, col_reg}<12'b101001100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101001100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101001100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101001100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101001100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101001100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b101001100101) && ({row_reg, col_reg}<12'b101001101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101001101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101001101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101001101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101001101011)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b101001101100) && ({row_reg, col_reg}<12'b101010000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101010000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101010001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b101010001001) && ({row_reg, col_reg}<12'b101010001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101010001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b101010001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b101010001101) && ({row_reg, col_reg}<12'b101010010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101010010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b101010010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101010010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101010010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b101010010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b101010010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b101010010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b101010010111) && ({row_reg, col_reg}<12'b101010011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101010011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101010011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101010011011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=12'b101010011100) && ({row_reg, col_reg}<12'b101010011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b101010011110) && ({row_reg, col_reg}<12'b101010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101010100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101010100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101010100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101010100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101010100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101010100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101010100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b101010100111) && ({row_reg, col_reg}<12'b101010101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101010101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101010101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b101010101100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=12'b101010101101) && ({row_reg, col_reg}<12'b101011000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101011000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101011001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101011001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101011001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101011001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101011001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101011001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101011001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101011001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b101011010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101011010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101011010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101011010011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b101011010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101011010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101011010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101011010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101011011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101011011001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101011011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b101011011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101011011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101011011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101011011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b101011011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101011100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101011100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101011100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101011100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b101011100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101011100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101011100110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b101011100111) && ({row_reg, col_reg}<12'b101100001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101100001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101100001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101100001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101100001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101100001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101100001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101100001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101100001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b101100010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101100010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b101100010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101100010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101100010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101100010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101100010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101100010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101100011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b101100011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101100011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101100011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101100011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101100011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101100011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101100011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101100100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101100100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101100100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101100100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101100100100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101100100101)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=12'b101100100110) && ({row_reg, col_reg}<12'b101101001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101101001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101101001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101101001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101101001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101101001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b101101001110) && ({row_reg, col_reg}<12'b101101010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101101010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101101010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b101101010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b101101010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101101010110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b101101010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101101011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101101011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101101011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b101101011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101101011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101101011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b101101011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101101011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101101100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101101100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b101101100010) && ({row_reg, col_reg}<12'b101101100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101101100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101101100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b101101100110) && ({row_reg, col_reg}<12'b101101101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101101101110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b101101101111) && ({row_reg, col_reg}<12'b101110000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101110000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b101110000011) && ({row_reg, col_reg}<12'b101110001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101110001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101110001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101110001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b101110001101) && ({row_reg, col_reg}<12'b101110001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101110001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b101110010000) && ({row_reg, col_reg}<12'b101110010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101110010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101110010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101110010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101110010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b101110010111) && ({row_reg, col_reg}<12'b101110011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101110011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b101110011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101110011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101110011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b101110011101) && ({row_reg, col_reg}<12'b101110100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101110100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101110100100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=12'b101110100101) && ({row_reg, col_reg}<12'b101111001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101111001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==12'b101111001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b101111001101) && ({row_reg, col_reg}<12'b101111010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b101111010101) && ({row_reg, col_reg}<12'b101111010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b101111010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101111011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b101111011001) && ({row_reg, col_reg}<12'b101111100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b101111100010) && ({row_reg, col_reg}<12'b101111100100)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=12'b101111100100) && ({row_reg, col_reg}<12'b110000010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b110000010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=12'b110000010010) && ({row_reg, col_reg}<12'b110000010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b110000010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b110000010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==12'b110000010111)) color_data = 12'b111011101110;



		if(({row_reg, col_reg}>=12'b110000011000) && ({row_reg, col_reg}<=12'b110010110010)) color_data = 12'b111111111111;
	end
endmodule