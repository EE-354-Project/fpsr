module steve_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}==10'b0000000000)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=10'b0000000001) && ({row_reg, col_reg}<10'b0000000100)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}>=10'b0000000100) && ({row_reg, col_reg}<10'b0000000111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0000000111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==10'b0000001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=10'b0000001001) && ({row_reg, col_reg}<10'b0000001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=10'b0000001100) && ({row_reg, col_reg}<10'b0000011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0000011000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=10'b0000011001) && ({row_reg, col_reg}<10'b0000011111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==10'b0000011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==10'b0000100000)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=10'b0000100001) && ({row_reg, col_reg}<10'b0000100111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0000100111)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==10'b0000101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0000101001)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==10'b0000101010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=10'b0000101011) && ({row_reg, col_reg}<10'b0000111000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0000111000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=10'b0000111001) && ({row_reg, col_reg}<10'b0000111111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==10'b0000111111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=10'b0001000000) && ({row_reg, col_reg}<10'b0001000010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=10'b0001000010) && ({row_reg, col_reg}<10'b0001000100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==10'b0001000100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==10'b0001000101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=10'b0001000110) && ({row_reg, col_reg}<10'b0001001000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=10'b0001001000) && ({row_reg, col_reg}<10'b0001001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==10'b0001001100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=10'b0001001101) && ({row_reg, col_reg}<10'b0001011000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=10'b0001011000) && ({row_reg, col_reg}<10'b0001011010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==10'b0001011010)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==10'b0001011011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=10'b0001011100) && ({row_reg, col_reg}<10'b0001011110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==10'b0001011110)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==10'b0001011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=10'b0001100000) && ({row_reg, col_reg}<10'b0001100100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=10'b0001100100) && ({row_reg, col_reg}<10'b0001101000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0001101000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=10'b0001101001) && ({row_reg, col_reg}<10'b0001101100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=10'b0001101100) && ({row_reg, col_reg}<10'b0001111111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==10'b0001111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=10'b0010000000) && ({row_reg, col_reg}<10'b0010001011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0010001011)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==10'b0010001100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==10'b0010001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==10'b0010001110)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=10'b0010001111) && ({row_reg, col_reg}<10'b0010011000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==10'b0010011000)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==10'b0010011001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0010011010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=10'b0010011011) && ({row_reg, col_reg}<10'b0010011111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==10'b0010011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=10'b0010100000) && ({row_reg, col_reg}<10'b0010101100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=10'b0010101100) && ({row_reg, col_reg}<10'b0010110000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=10'b0010110000) && ({row_reg, col_reg}<10'b0010111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=10'b0010111000) && ({row_reg, col_reg}<10'b0010111011)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=10'b0010111011) && ({row_reg, col_reg}<10'b0010111111)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==10'b0010111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=10'b0011000000) && ({row_reg, col_reg}<10'b0011000010)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=10'b0011000010) && ({row_reg, col_reg}<10'b0011001000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0011001000)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=10'b0011001001) && ({row_reg, col_reg}<10'b0011001100)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=10'b0011001100) && ({row_reg, col_reg}<10'b0011010000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=10'b0011010000) && ({row_reg, col_reg}<10'b0011010100)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}>=10'b0011010100) && ({row_reg, col_reg}<10'b0011010110)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}>=10'b0011010110) && ({row_reg, col_reg}<10'b0011011000)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==10'b0011011000)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=10'b0011011001) && ({row_reg, col_reg}<10'b0011011110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0011011110)) color_data = 12'b000100010000;

		if(({row_reg, col_reg}==10'b0011011111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}>=10'b0011100000) && ({row_reg, col_reg}<10'b0011100100)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=10'b0011100100) && ({row_reg, col_reg}<10'b0011101000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==10'b0011101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=10'b0011101001) && ({row_reg, col_reg}<10'b0011101011)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}>=10'b0011101011) && ({row_reg, col_reg}<10'b0011110000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=10'b0011110000) && ({row_reg, col_reg}<10'b0011110011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}>=10'b0011110011) && ({row_reg, col_reg}<10'b0011110110)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=10'b0011110110) && ({row_reg, col_reg}<10'b0011111000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==10'b0011111000)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==10'b0011111001)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==10'b0011111010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=10'b0011111011) && ({row_reg, col_reg}<10'b0011111101)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==10'b0011111101)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==10'b0011111110)) color_data = 12'b001000010000;

		if(({row_reg, col_reg}==10'b0011111111)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==10'b0100000000)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}>=10'b0100000001) && ({row_reg, col_reg}<10'b0100000011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0100000011)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==10'b0100000100)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=10'b0100000101) && ({row_reg, col_reg}<10'b0100001000)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=10'b0100001000) && ({row_reg, col_reg}<10'b0100001101)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}>=10'b0100001101) && ({row_reg, col_reg}<10'b0100010000)) color_data = 12'b101110010111;
		if(({row_reg, col_reg}==10'b0100010000)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0100010001)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b0100010010)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0100010011)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b0100010100)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0100010101)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b0100010110)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0100010111)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b0100011000) && ({row_reg, col_reg}<10'b0100011010)) color_data = 12'b100101110101;
		if(({row_reg, col_reg}==10'b0100011010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==10'b0100011011)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==10'b0100011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=10'b0100011101) && ({row_reg, col_reg}<10'b0100011111)) color_data = 12'b001100100000;

		if(({row_reg, col_reg}==10'b0100011111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==10'b0100100000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0100100001)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==10'b0100100010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==10'b0100100011)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==10'b0100100100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=10'b0100100101) && ({row_reg, col_reg}<10'b0100101001)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}>=10'b0100101001) && ({row_reg, col_reg}<10'b0100101100)) color_data = 12'b110010000111;
		if(({row_reg, col_reg}>=10'b0100101100) && ({row_reg, col_reg}<10'b0100110000)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}>=10'b0100110000) && ({row_reg, col_reg}<10'b0100110010)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0100110010)) color_data = 12'b101110010111;
		if(({row_reg, col_reg}==10'b0100110011)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}>=10'b0100110100) && ({row_reg, col_reg}<10'b0100110110)) color_data = 12'b110010000111;
		if(({row_reg, col_reg}==10'b0100110110)) color_data = 12'b110010010111;
		if(({row_reg, col_reg}==10'b0100110111)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}>=10'b0100111000) && ({row_reg, col_reg}<10'b0100111011)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b0100111011)) color_data = 12'b100101110101;
		if(({row_reg, col_reg}==10'b0100111100)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==10'b0100111101)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==10'b0100111110)) color_data = 12'b001100010000;

		if(({row_reg, col_reg}==10'b0100111111)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==10'b0101000000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=10'b0101000001) && ({row_reg, col_reg}<10'b0101000011)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==10'b0101000011)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}>=10'b0101000100) && ({row_reg, col_reg}<10'b0101000111)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}>=10'b0101000111) && ({row_reg, col_reg}<10'b0101001100)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}>=10'b0101001100) && ({row_reg, col_reg}<10'b0101010000)) color_data = 12'b110010010111;
		if(({row_reg, col_reg}>=10'b0101010000) && ({row_reg, col_reg}<10'b0101010011)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0101010011)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b0101010100)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0101010101)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b0101010110)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0101010111)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b0101011000)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}>=10'b0101011001) && ({row_reg, col_reg}<10'b0101011100)) color_data = 12'b100101110101;
		if(({row_reg, col_reg}>=10'b0101011100) && ({row_reg, col_reg}<10'b0101011110)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==10'b0101011110)) color_data = 12'b001100100000;

		if(({row_reg, col_reg}==10'b0101011111)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==10'b0101100000)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}>=10'b0101100001) && ({row_reg, col_reg}<10'b0101100011)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==10'b0101100011)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==10'b0101100100)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b0101100101)) color_data = 12'b101110010111;
		if(({row_reg, col_reg}==10'b0101100110)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0101100111)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b0101101000) && ({row_reg, col_reg}<10'b0101101100)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}>=10'b0101101100) && ({row_reg, col_reg}<10'b0101110000)) color_data = 12'b110010010111;
		if(({row_reg, col_reg}>=10'b0101110000) && ({row_reg, col_reg}<10'b0101110011)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0101110011)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b0101110100) && ({row_reg, col_reg}<10'b0101110111)) color_data = 12'b110010010111;
		if(({row_reg, col_reg}==10'b0101110111)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}>=10'b0101111000) && ({row_reg, col_reg}<10'b0101111010)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}==10'b0101111010)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b0101111011)) color_data = 12'b100101110101;
		if(({row_reg, col_reg}==10'b0101111100)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==10'b0101111101)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}==10'b0101111110)) color_data = 12'b010000100000;

		if(({row_reg, col_reg}==10'b0101111111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==10'b0110000000)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==10'b0110000001)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b0110000010)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b0110000011)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b0110000100)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0110000101)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}>=10'b0110000110) && ({row_reg, col_reg}<10'b0110001000)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b0110001000) && ({row_reg, col_reg}<10'b0110001100)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}>=10'b0110001100) && ({row_reg, col_reg}<10'b0110001110)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b0110001110) && ({row_reg, col_reg}<10'b0110010000)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}>=10'b0110010000) && ({row_reg, col_reg}<10'b0110010100)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}==10'b0110010100)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b0110010101)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}>=10'b0110010110) && ({row_reg, col_reg}<10'b0110011000)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b0110011000)) color_data = 12'b101001100101;
		if(({row_reg, col_reg}>=10'b0110011001) && ({row_reg, col_reg}<10'b0110011101)) color_data = 12'b100101100100;

		if(({row_reg, col_reg}>=10'b0110011101) && ({row_reg, col_reg}<10'b0110100000)) color_data = 12'b100101100101;
		if(({row_reg, col_reg}>=10'b0110100000) && ({row_reg, col_reg}<10'b0110100100)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b0110100100)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b0110100101) && ({row_reg, col_reg}<10'b0110100111)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0110100111)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b0110101000)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b0110101001)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}>=10'b0110101010) && ({row_reg, col_reg}<10'b0110101100)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}>=10'b0110101100) && ({row_reg, col_reg}<10'b0110101110)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}>=10'b0110101110) && ({row_reg, col_reg}<10'b0110110000)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}>=10'b0110110000) && ({row_reg, col_reg}<10'b0110110010)) color_data = 12'b100101100101;
		if(({row_reg, col_reg}==10'b0110110010)) color_data = 12'b101001100101;
		if(({row_reg, col_reg}==10'b0110110011)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}==10'b0110110100)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}>=10'b0110110101) && ({row_reg, col_reg}<10'b0110110111)) color_data = 12'b110010000111;
		if(({row_reg, col_reg}==10'b0110110111)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b0110111000) && ({row_reg, col_reg}<10'b0110111010)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==10'b0110111010)) color_data = 12'b101001100101;
		if(({row_reg, col_reg}>=10'b0110111011) && ({row_reg, col_reg}<10'b0110111111)) color_data = 12'b100101100100;

		if(({row_reg, col_reg}==10'b0110111111)) color_data = 12'b100101100101;
		if(({row_reg, col_reg}>=10'b0111000000) && ({row_reg, col_reg}<10'b0111000100)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}>=10'b0111000100) && ({row_reg, col_reg}<10'b0111000110)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b0111000110)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b0111000111)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b0111001000)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b0111001001)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}>=10'b0111001010) && ({row_reg, col_reg}<10'b0111001100)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}>=10'b0111001100) && ({row_reg, col_reg}<10'b0111010000)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}>=10'b0111010000) && ({row_reg, col_reg}<10'b0111010010)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}>=10'b0111010010) && ({row_reg, col_reg}<10'b0111010100)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}>=10'b0111010100) && ({row_reg, col_reg}<10'b0111010111)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b0111010111)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b0111011000) && ({row_reg, col_reg}<10'b0111011111)) color_data = 12'b100101100100;

		if(({row_reg, col_reg}==10'b0111011111)) color_data = 12'b100101100101;
		if(({row_reg, col_reg}>=10'b0111100000) && ({row_reg, col_reg}<10'b0111100010)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b0111100010)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b0111100011)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b0111100100)) color_data = 12'b101110010111;
		if(({row_reg, col_reg}==10'b0111100101)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==10'b0111100110)) color_data = 12'b101110010111;
		if(({row_reg, col_reg}==10'b0111100111)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}>=10'b0111101000) && ({row_reg, col_reg}<10'b0111101100)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==10'b0111101100)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b0111101101)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b0111101110)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b0111101111)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b0111110000)) color_data = 12'b100101100101;
		if(({row_reg, col_reg}==10'b0111110001)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}==10'b0111110010)) color_data = 12'b100101110101;
		if(({row_reg, col_reg}==10'b0111110011)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=10'b0111110100) && ({row_reg, col_reg}<10'b0111110111)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==10'b0111110111)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==10'b0111111000)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==10'b0111111001)) color_data = 12'b100101110101;
		if(({row_reg, col_reg}==10'b0111111010)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==10'b0111111011)) color_data = 12'b101001110110;

		if(({row_reg, col_reg}>=10'b0111111100) && ({row_reg, col_reg}<10'b1000000000)) color_data = 12'b100101100101;
		if(({row_reg, col_reg}==10'b1000000000)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b1000000001)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1000000010)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b1000000011)) color_data = 12'b101110010111;
		if(({row_reg, col_reg}==10'b1000000100)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==10'b1000000101)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==10'b1000000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==10'b1000000111)) color_data = 12'b111111101110;
		if(({row_reg, col_reg}==10'b1000001000)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}>=10'b1000001001) && ({row_reg, col_reg}<10'b1000001011)) color_data = 12'b010100110111;
		if(({row_reg, col_reg}==10'b1000001011)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==10'b1000001100)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b1000001101)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b1000001110) && ({row_reg, col_reg}<10'b1000010000)) color_data = 12'b101101110101;
		if(({row_reg, col_reg}>=10'b1000010000) && ({row_reg, col_reg}<10'b1000010010)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b1000010010)) color_data = 12'b101110010111;
		if(({row_reg, col_reg}==10'b1000010011)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==10'b1000010100)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==10'b1000010101)) color_data = 12'b010100110111;
		if(({row_reg, col_reg}==10'b1000010110)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==10'b1000010111)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==10'b1000011000)) color_data = 12'b111111101110;
		if(({row_reg, col_reg}>=10'b1000011001) && ({row_reg, col_reg}<10'b1000011011)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==10'b1000011011)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==10'b1000011100)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}>=10'b1000011101) && ({row_reg, col_reg}<10'b1000011111)) color_data = 12'b101001110110;

		if(({row_reg, col_reg}==10'b1000011111)) color_data = 12'b101001110111;
		if(({row_reg, col_reg}==10'b1000100000)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b1000100001)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1000100010)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b1000100011)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==10'b1000100100)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}>=10'b1000100101) && ({row_reg, col_reg}<10'b1000100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==10'b1000100111)) color_data = 12'b111111101111;
		if(({row_reg, col_reg}==10'b1000101000)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==10'b1000101001)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==10'b1000101010)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==10'b1000101011)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==10'b1000101100)) color_data = 12'b101001110111;
		if(({row_reg, col_reg}==10'b1000101101)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b1000101110)) color_data = 12'b101101110101;
		if(({row_reg, col_reg}==10'b1000101111)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}==10'b1000110000)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1000110001)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b1000110010)) color_data = 12'b101110010111;
		if(({row_reg, col_reg}==10'b1000110011)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==10'b1000110100)) color_data = 12'b010100110111;
		if(({row_reg, col_reg}==10'b1000110101)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==10'b1000110110)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==10'b1000110111)) color_data = 12'b010101011000;
		if(({row_reg, col_reg}>=10'b1000111000) && ({row_reg, col_reg}<10'b1000111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==10'b1000111011)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}>=10'b1000111100) && ({row_reg, col_reg}<10'b1000111110)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b1000111110)) color_data = 12'b101001110110;

		if(({row_reg, col_reg}==10'b1000111111)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==10'b1001000000)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}>=10'b1001000001) && ({row_reg, col_reg}<10'b1001000100)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}>=10'b1001000100) && ({row_reg, col_reg}<10'b1001000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==10'b1001000111)) color_data = 12'b111111101111;
		if(({row_reg, col_reg}==10'b1001001000)) color_data = 12'b010101000111;
		if(({row_reg, col_reg}>=10'b1001001001) && ({row_reg, col_reg}<10'b1001001011)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==10'b1001001011)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==10'b1001001100)) color_data = 12'b101001110111;
		if(({row_reg, col_reg}>=10'b1001001101) && ({row_reg, col_reg}<10'b1001001111)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b1001001111)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}==10'b1001010000)) color_data = 12'b110010000111;
		if(({row_reg, col_reg}>=10'b1001010001) && ({row_reg, col_reg}<10'b1001010011)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1001010011)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==10'b1001010100)) color_data = 12'b011000110111;
		if(({row_reg, col_reg}==10'b1001010101)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==10'b1001010110)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==10'b1001010111)) color_data = 12'b010101011000;
		if(({row_reg, col_reg}>=10'b1001011000) && ({row_reg, col_reg}<10'b1001011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==10'b1001011011)) color_data = 12'b111111101110;
		if(({row_reg, col_reg}==10'b1001011100)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=10'b1001011101) && ({row_reg, col_reg}<10'b1001011111)) color_data = 12'b101001110110;

		if(({row_reg, col_reg}==10'b1001011111)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}>=10'b1001100000) && ({row_reg, col_reg}<10'b1001100010)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b1001100010)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b1001100011)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1001100100)) color_data = 12'b111111101110;
		if(({row_reg, col_reg}==10'b1001100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==10'b1001100110)) color_data = 12'b111111101111;
		if(({row_reg, col_reg}==10'b1001100111)) color_data = 12'b111111011110;
		if(({row_reg, col_reg}==10'b1001101000)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==10'b1001101001)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==10'b1001101010)) color_data = 12'b010100110111;
		if(({row_reg, col_reg}==10'b1001101011)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==10'b1001101100)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==10'b1001101101)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b1001101110) && ({row_reg, col_reg}<10'b1001110000)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b1001110000)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}>=10'b1001110001) && ({row_reg, col_reg}<10'b1001110011)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1001110011)) color_data = 12'b101001110111;
		if(({row_reg, col_reg}==10'b1001110100)) color_data = 12'b011101000110;
		if(({row_reg, col_reg}==10'b1001110101)) color_data = 12'b010100110111;
		if(({row_reg, col_reg}==10'b1001110110)) color_data = 12'b010101000111;
		if(({row_reg, col_reg}==10'b1001110111)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==10'b1001111000)) color_data = 12'b111111101110;
		if(({row_reg, col_reg}>=10'b1001111001) && ({row_reg, col_reg}<10'b1001111011)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==10'b1001111011)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==10'b1001111100)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}>=10'b1001111101) && ({row_reg, col_reg}<10'b1001111111)) color_data = 12'b101001110101;

		if(({row_reg, col_reg}==10'b1001111111)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b1010000000)) color_data = 12'b100101010011;
		if(({row_reg, col_reg}>=10'b1010000001) && ({row_reg, col_reg}<10'b1010000011)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}==10'b1010000011)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}>=10'b1010000100) && ({row_reg, col_reg}<10'b1010000111)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}>=10'b1010000111) && ({row_reg, col_reg}<10'b1010001001)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==10'b1010001001)) color_data = 12'b101001111000;
		if(({row_reg, col_reg}==10'b1010001010)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==10'b1010001011)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==10'b1010001100)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=10'b1010001101) && ({row_reg, col_reg}<10'b1010001111)) color_data = 12'b011100110010;
		if(({row_reg, col_reg}==10'b1010001111)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1010010000)) color_data = 12'b011101000100;
		if(({row_reg, col_reg}>=10'b1010010001) && ({row_reg, col_reg}<10'b1010010011)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==10'b1010010011)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1010010100)) color_data = 12'b101001110111;
		if(({row_reg, col_reg}==10'b1010010101)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}==10'b1010010110)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==10'b1010010111)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}>=10'b1010011000) && ({row_reg, col_reg}<10'b1010011010)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}>=10'b1010011010) && ({row_reg, col_reg}<10'b1010011100)) color_data = 12'b100101110101;
		if(({row_reg, col_reg}>=10'b1010011100) && ({row_reg, col_reg}<10'b1010011110)) color_data = 12'b100001010011;

		if(({row_reg, col_reg}>=10'b1010011110) && ({row_reg, col_reg}<10'b1010100000)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==10'b1010100000)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}==10'b1010100001)) color_data = 12'b101001010011;
		if(({row_reg, col_reg}==10'b1010100010)) color_data = 12'b101001010100;
		if(({row_reg, col_reg}==10'b1010100011)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}==10'b1010100100)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}==10'b1010100101)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b1010100110)) color_data = 12'b101110000101;
		if(({row_reg, col_reg}==10'b1010100111)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}==10'b1010101000)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1010101001)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b1010101010)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1010101011)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}>=10'b1010101100) && ({row_reg, col_reg}<10'b1010101110)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==10'b1010101110)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}>=10'b1010101111) && ({row_reg, col_reg}<10'b1010110001)) color_data = 12'b011000110011;
		if(({row_reg, col_reg}==10'b1010110001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=10'b1010110010) && ({row_reg, col_reg}<10'b1010110100)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==10'b1010110100)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1010110101)) color_data = 12'b110010000111;
		if(({row_reg, col_reg}==10'b1010110110)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1010110111)) color_data = 12'b110010000110;
		if(({row_reg, col_reg}==10'b1010111000)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==10'b1010111001)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}>=10'b1010111010) && ({row_reg, col_reg}<10'b1010111100)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==10'b1010111100)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==10'b1010111101)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==10'b1010111110)) color_data = 12'b011101010010;

		if(({row_reg, col_reg}==10'b1010111111)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==10'b1011000000)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}>=10'b1011000001) && ({row_reg, col_reg}<10'b1011000011)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==10'b1011000011)) color_data = 12'b101001100101;
		if(({row_reg, col_reg}>=10'b1011000100) && ({row_reg, col_reg}<10'b1011000110)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b1011000110)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}==10'b1011000111)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}>=10'b1011001000) && ({row_reg, col_reg}<10'b1011001011)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1011001011)) color_data = 12'b101010000110;
		if(({row_reg, col_reg}==10'b1011001100)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==10'b1011001101)) color_data = 12'b011000110010;
		if(({row_reg, col_reg}>=10'b1011001110) && ({row_reg, col_reg}<10'b1011010001)) color_data = 12'b011000110011;
		if(({row_reg, col_reg}==10'b1011010001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==10'b1011010010)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==10'b1011010011)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==10'b1011010100)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}>=10'b1011010101) && ({row_reg, col_reg}<10'b1011011000)) color_data = 12'b110010000110;
		if(({row_reg, col_reg}==10'b1011011000)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}==10'b1011011001)) color_data = 12'b101001110100;
		if(({row_reg, col_reg}==10'b1011011010)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}==10'b1011011011)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==10'b1011011100)) color_data = 12'b100001010011;

		if(({row_reg, col_reg}>=10'b1011011101) && ({row_reg, col_reg}<10'b1011100000)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}>=10'b1011100000) && ({row_reg, col_reg}<10'b1011100100)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}>=10'b1011100100) && ({row_reg, col_reg}<10'b1011100110)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}==10'b1011100110)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b1011100111)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}>=10'b1011101000) && ({row_reg, col_reg}<10'b1011101010)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b1011101010)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==10'b1011101011)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==10'b1011101100)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1011101101)) color_data = 12'b011000110010;
		if(({row_reg, col_reg}>=10'b1011101110) && ({row_reg, col_reg}<10'b1011110000)) color_data = 12'b011000110011;
		if(({row_reg, col_reg}==10'b1011110000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==10'b1011110001)) color_data = 12'b011000110011;
		if(({row_reg, col_reg}==10'b1011110010)) color_data = 12'b011000110010;
		if(({row_reg, col_reg}==10'b1011110011)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==10'b1011110100)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}>=10'b1011110101) && ({row_reg, col_reg}<10'b1011110111)) color_data = 12'b101110000110;
		if(({row_reg, col_reg}==10'b1011110111)) color_data = 12'b101101110101;
		if(({row_reg, col_reg}>=10'b1011111000) && ({row_reg, col_reg}<10'b1011111010)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}>=10'b1011111010) && ({row_reg, col_reg}<10'b1011111100)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==10'b1011111100)) color_data = 12'b100001000011;

		if(({row_reg, col_reg}>=10'b1011111101) && ({row_reg, col_reg}<10'b1100000001)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==10'b1100000001)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}>=10'b1100000010) && ({row_reg, col_reg}<10'b1100000101)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}>=10'b1100000101) && ({row_reg, col_reg}<10'b1100000111)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==10'b1100000111)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}>=10'b1100001000) && ({row_reg, col_reg}<10'b1100011000)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1100011000)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==10'b1100011001)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}>=10'b1100011010) && ({row_reg, col_reg}<10'b1100011100)) color_data = 12'b100101010100;

		if(({row_reg, col_reg}>=10'b1100011100) && ({row_reg, col_reg}<10'b1100100001)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1100100001) && ({row_reg, col_reg}<10'b1100100100)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}>=10'b1100100100) && ({row_reg, col_reg}<10'b1100101000)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}>=10'b1100101000) && ({row_reg, col_reg}<10'b1100101010)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1100101010)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}>=10'b1100101011) && ({row_reg, col_reg}<10'b1100110000)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1100110000)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}>=10'b1100110001) && ({row_reg, col_reg}<10'b1100110011)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1100110011)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}==10'b1100110100)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1100110101)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}>=10'b1100110110) && ({row_reg, col_reg}<10'b1100111000)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=10'b1100111000) && ({row_reg, col_reg}<10'b1100111100)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}>=10'b1100111100) && ({row_reg, col_reg}<10'b1100111111)) color_data = 12'b100001000011;

		if(({row_reg, col_reg}==10'b1100111111)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1101000000) && ({row_reg, col_reg}<10'b1101000010)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==10'b1101000010)) color_data = 12'b100001100100;
		if(({row_reg, col_reg}>=10'b1101000011) && ({row_reg, col_reg}<10'b1101000101)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}==10'b1101000101)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}>=10'b1101000110) && ({row_reg, col_reg}<10'b1101001000)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}>=10'b1101001000) && ({row_reg, col_reg}<10'b1101001010)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=10'b1101001010) && ({row_reg, col_reg}<10'b1101001100)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}>=10'b1101001100) && ({row_reg, col_reg}<10'b1101011000)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1101011000)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==10'b1101011001)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==10'b1101011010)) color_data = 12'b100101010011;
		if(({row_reg, col_reg}==10'b1101011011)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}>=10'b1101011100) && ({row_reg, col_reg}<10'b1101011111)) color_data = 12'b100001010011;

		if(({row_reg, col_reg}>=10'b1101011111) && ({row_reg, col_reg}<10'b1101100101)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}>=10'b1101100101) && ({row_reg, col_reg}<10'b1101101000)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}>=10'b1101101000) && ({row_reg, col_reg}<10'b1101110000)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1101110000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=10'b1101110001) && ({row_reg, col_reg}<10'b1101111000)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=10'b1101111000) && ({row_reg, col_reg}<10'b1101111101)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1101111101) && ({row_reg, col_reg}<10'b1101111111)) color_data = 12'b011101010011;

		if(({row_reg, col_reg}==10'b1101111111)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==10'b1110000000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=10'b1110000001) && ({row_reg, col_reg}<10'b1110000100)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=10'b1110000100) && ({row_reg, col_reg}<10'b1110000111)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==10'b1110000111)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=10'b1110001000) && ({row_reg, col_reg}<10'b1110001010)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}>=10'b1110001010) && ({row_reg, col_reg}<10'b1110001100)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}>=10'b1110001100) && ({row_reg, col_reg}<10'b1110001111)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==10'b1110001111)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1110010000) && ({row_reg, col_reg}<10'b1110010100)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=10'b1110010100) && ({row_reg, col_reg}<10'b1110010110)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==10'b1110010110)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=10'b1110010111) && ({row_reg, col_reg}<10'b1110011100)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1110011100) && ({row_reg, col_reg}<10'b1110011111)) color_data = 12'b011101000011;

		if(({row_reg, col_reg}==10'b1110011111)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==10'b1110100000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=10'b1110100001) && ({row_reg, col_reg}<10'b1110100100)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=10'b1110100100) && ({row_reg, col_reg}<10'b1110100110)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=10'b1110100110) && ({row_reg, col_reg}<10'b1110101000)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==10'b1110101000)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}>=10'b1110101001) && ({row_reg, col_reg}<10'b1110101011)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}>=10'b1110101011) && ({row_reg, col_reg}<10'b1110101101)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==10'b1110101101)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}>=10'b1110101110) && ({row_reg, col_reg}<10'b1110110000)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1110110000) && ({row_reg, col_reg}<10'b1110110100)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=10'b1110110100) && ({row_reg, col_reg}<10'b1110110110)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}>=10'b1110110110) && ({row_reg, col_reg}<10'b1110111100)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1110111100) && ({row_reg, col_reg}<10'b1110111111)) color_data = 12'b011101000011;

		if(({row_reg, col_reg}==10'b1110111111)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==10'b1111000000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=10'b1111000001) && ({row_reg, col_reg}<10'b1111000100)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=10'b1111000100) && ({row_reg, col_reg}<10'b1111000110)) color_data = 12'b011100110010;
		if(({row_reg, col_reg}>=10'b1111000110) && ({row_reg, col_reg}<10'b1111001000)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}>=10'b1111001000) && ({row_reg, col_reg}<10'b1111001010)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==10'b1111001010)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==10'b1111001011)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1111001100) && ({row_reg, col_reg}<10'b1111001110)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==10'b1111001110)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1111001111)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}>=10'b1111010000) && ({row_reg, col_reg}<10'b1111010100)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=10'b1111010100) && ({row_reg, col_reg}<10'b1111011010)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==10'b1111011010)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==10'b1111011011)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1111011100) && ({row_reg, col_reg}<10'b1111011110)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==10'b1111011110)) color_data = 12'b011101000011;

		if(({row_reg, col_reg}==10'b1111011111)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}>=10'b1111100000) && ({row_reg, col_reg}<10'b1111100010)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==10'b1111100010)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=10'b1111100011) && ({row_reg, col_reg}<10'b1111100110)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=10'b1111100110) && ({row_reg, col_reg}<10'b1111101000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=10'b1111101000) && ({row_reg, col_reg}<10'b1111101101)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1111101101) && ({row_reg, col_reg}<10'b1111110000)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==10'b1111110000)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1111110001) && ({row_reg, col_reg}<10'b1111110011)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==10'b1111110011)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1111110100) && ({row_reg, col_reg}<10'b1111110110)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}>=10'b1111110110) && ({row_reg, col_reg}<10'b1111111001)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=10'b1111111001) && ({row_reg, col_reg}<10'b1111111100)) color_data = 12'b100001010100;

		if(({row_reg, col_reg}>=10'b1111111100) && ({row_reg, col_reg}<=10'b1111111111)) color_data = 12'b011101010011;
	end
endmodule