module g1_rom (
    input wire clk,
    input wire [3:0] row,
    input wire [6:0] col,
    output reg [11:0] color_data
);

    (* rom_style = "block" *)

    reg [3:0] row_reg;
    reg [6:0] col_reg;

    always @(posedge clk) begin
        row_reg <= row;
        col_reg <= col;
    end

    always @(*) begin
        case ({row_reg, col_reg})
            11'b00000000000: color_data = 12'b111111111111;
            11'b00000000001: color_data = 12'b111111111111;
            11'b00000000010: color_data = 12'b111111111111;
            11'b00000000011: color_data = 12'b111111111111;
            11'b00000000100: color_data = 12'b111111111111;
            11'b00000000101: color_data = 12'b111111111111;
            11'b00000000110: color_data = 12'b111111111111;
            11'b00000000111: color_data = 12'b111111111111;
            11'b00000001000: color_data = 12'b111111111111;
            11'b00000001001: color_data = 12'b111111111111;
            11'b00000001010: color_data = 12'b111111111111;
            11'b00000001011: color_data = 12'b111111111111;
            11'b00000001100: color_data = 12'b111111111111;
            11'b00000001101: color_data = 12'b111111111111;
            11'b00000001110: color_data = 12'b111111111111;
            11'b00000001111: color_data = 12'b111111111111;
            11'b00000010000: color_data = 12'b111111111111;
            11'b00000010001: color_data = 12'b111111111111;
            11'b00000010010: color_data = 12'b111111111111;
            11'b00000010011: color_data = 12'b111111111111;
            11'b00000010100: color_data = 12'b111111111111;
            11'b00000010101: color_data = 12'b111111111111;
            11'b00000010110: color_data = 12'b111111111111;
            11'b00000010111: color_data = 12'b111111111111;
            11'b00000011000: color_data = 12'b111111111111;
            11'b00000011001: color_data = 12'b111111111111;
            11'b00000011010: color_data = 12'b111111111111;
            11'b00000011011: color_data = 12'b111111111111;
            11'b00000011100: color_data = 12'b111111111111;
            11'b00000011101: color_data = 12'b111111111111;
            11'b00000011110: color_data = 12'b111111111111;
            11'b00000011111: color_data = 12'b111111111111;
            11'b00000100000: color_data = 12'b111111111111;
            11'b00000100001: color_data = 12'b111111111111;
            11'b00000100010: color_data = 12'b111111111111;
            11'b00000100011: color_data = 12'b111111111111;
            11'b00000100100: color_data = 12'b111111111111;
            11'b00000100101: color_data = 12'b111111111111;
            11'b00000100110: color_data = 12'b111111111111;
            11'b00000100111: color_data = 12'b111111111111;
            11'b00000101000: color_data = 12'b111111111111;
            11'b00000101001: color_data = 12'b111111111111;
            11'b00000101010: color_data = 12'b111111111111;
            11'b00000101011: color_data = 12'b111111111111;
            11'b00000101100: color_data = 12'b111111111111;
            11'b00000101101: color_data = 12'b111111111111;
            11'b00000101110: color_data = 12'b111111111111;
            11'b00000101111: color_data = 12'b111111111111;
            11'b00000110000: color_data = 12'b111111111111;
            11'b00000110001: color_data = 12'b111111111111;
            11'b00000110010: color_data = 12'b111111111111;
            11'b00000110011: color_data = 12'b111111111111;
            11'b00000110100: color_data = 12'b111111111111;
            11'b00000110101: color_data = 12'b111111111111;
            11'b00000110110: color_data = 12'b111111111111;
            11'b00000110111: color_data = 12'b111111111111;
            11'b00000111000: color_data = 12'b111111111111;
            11'b00000111001: color_data = 12'b111111111111;
            11'b00000111010: color_data = 12'b111111111111;
            11'b00000111011: color_data = 12'b111111111111;
            11'b00000111100: color_data = 12'b111111111111;
            11'b00000111101: color_data = 12'b111111111111;
            11'b00000111110: color_data = 12'b111111111111;
            11'b00000111111: color_data = 12'b111111111111;
            11'b00001000000: color_data = 12'b111111111111;
            11'b00001000001: color_data = 12'b111111111111;
            11'b00001000010: color_data = 12'b111111111111;
            11'b00001000011: color_data = 12'b111111111111;
            11'b00001000100: color_data = 12'b111111111111;
            11'b00001000101: color_data = 12'b111111111111;
            11'b00001000110: color_data = 12'b111111111111;
            11'b00001000111: color_data = 12'b111111111111;
            11'b00001001000: color_data = 12'b111111111111;
            11'b00001001001: color_data = 12'b111111111111;
            11'b00001001010: color_data = 12'b111111111111;
            11'b00001001011: color_data = 12'b111111111111;
            11'b00001001100: color_data = 12'b111111111111;
            11'b00001001101: color_data = 12'b111111111111;
            11'b00010000000: color_data = 12'b111111111111;
            11'b00010000001: color_data = 12'b111111111111;
            11'b00010000010: color_data = 12'b111111111111;
            11'b00010000011: color_data = 12'b111111111111;
            11'b00010000100: color_data = 12'b111111111111;
            11'b00010000101: color_data = 12'b111111111111;
            11'b00010000110: color_data = 12'b111111111111;
            11'b00010000111: color_data = 12'b111111111111;
            11'b00010001000: color_data = 12'b111111111111;
            11'b00010001001: color_data = 12'b111111111111;
            11'b00010001010: color_data = 12'b111111111111;
            11'b00010001011: color_data = 12'b111111111111;
            11'b00010001100: color_data = 12'b111111111111;
            11'b00010001101: color_data = 12'b111111111111;
            11'b00010001110: color_data = 12'b111111111111;
            11'b00010001111: color_data = 12'b111111111111;
            11'b00010010000: color_data = 12'b111111111111;
            11'b00010010001: color_data = 12'b111111111111;
            11'b00010010010: color_data = 12'b111111111111;
            11'b00010010011: color_data = 12'b111111111111;
            11'b00010010100: color_data = 12'b111111111111;
            11'b00010010101: color_data = 12'b111111111111;
            11'b00010010110: color_data = 12'b111111111111;
            11'b00010010111: color_data = 12'b111111111111;
            11'b00010011000: color_data = 12'b111111111111;
            11'b00010011001: color_data = 12'b111111111111;
            11'b00010011010: color_data = 12'b111111111111;
            11'b00010011011: color_data = 12'b111111111111;
            11'b00010011100: color_data = 12'b111111111111;
            11'b00010011101: color_data = 12'b111111111111;
            11'b00010011110: color_data = 12'b111111111111;
            11'b00010011111: color_data = 12'b111111111111;
            11'b00010100000: color_data = 12'b111111111111;
            11'b00010100001: color_data = 12'b111111111111;
            11'b00010100010: color_data = 12'b111111111111;
            11'b00010100011: color_data = 12'b111111111111;
            11'b00010100100: color_data = 12'b111111111111;
            11'b00010100101: color_data = 12'b111111111111;
            11'b00010100110: color_data = 12'b111111111111;
            11'b00010100111: color_data = 12'b111111111111;
            11'b00010101000: color_data = 12'b111111111111;
            11'b00010101001: color_data = 12'b111111111111;
            11'b00010101010: color_data = 12'b111111111111;
            11'b00010101011: color_data = 12'b111111111111;
            11'b00010101100: color_data = 12'b111111111111;
            11'b00010101101: color_data = 12'b111111111111;
            11'b00010101110: color_data = 12'b111111111111;
            11'b00010101111: color_data = 12'b111111111111;
            11'b00010110000: color_data = 12'b111111111111;
            11'b00010110001: color_data = 12'b111111111111;
            11'b00010110010: color_data = 12'b111111111111;
            11'b00010110011: color_data = 12'b111111111111;
            11'b00010110100: color_data = 12'b111111111111;
            11'b00010110101: color_data = 12'b111111111111;
            11'b00010110110: color_data = 12'b111111111111;
            11'b00010110111: color_data = 12'b111111111111;
            11'b00010111000: color_data = 12'b111111111111;
            11'b00010111001: color_data = 12'b111111111111;
            11'b00010111010: color_data = 12'b111111111111;
            11'b00010111011: color_data = 12'b111111111111;
            11'b00010111100: color_data = 12'b111111111111;
            11'b00010111101: color_data = 12'b111111111111;
            11'b00010111110: color_data = 12'b111111111111;
            11'b00010111111: color_data = 12'b111111111111;
            11'b00011000000: color_data = 12'b111111111111;
            11'b00011000001: color_data = 12'b111111111111;
            11'b00011000010: color_data = 12'b111111111111;
            11'b00011000011: color_data = 12'b111111111111;
            11'b00011000100: color_data = 12'b111111111111;
            11'b00011000101: color_data = 12'b111111111111;
            11'b00011000110: color_data = 12'b111111111111;
            11'b00011000111: color_data = 12'b111111111111;
            11'b00011001000: color_data = 12'b111111111111;
            11'b00011001001: color_data = 12'b111111111111;
            11'b00011001010: color_data = 12'b111111111111;
            11'b00011001011: color_data = 12'b111111111111;
            11'b00011001100: color_data = 12'b111111111111;
            11'b00011001101: color_data = 12'b111111111111;
            11'b00100000000: color_data = 12'b111111111111;
            11'b00100000001: color_data = 12'b111111111111;
            11'b00100000010: color_data = 12'b111111111111;
            11'b00100000011: color_data = 12'b111111111111;
            11'b00100000100: color_data = 12'b111111111111;
            11'b00100000101: color_data = 12'b111111111111;
            11'b00100000110: color_data = 12'b111111111111;
            11'b00100000111: color_data = 12'b111111111111;
            11'b00100001000: color_data = 12'b111111111111;
            11'b00100001001: color_data = 12'b111111111111;
            11'b00100001010: color_data = 12'b111111111111;
            11'b00100001011: color_data = 12'b111111111111;
            11'b00100001100: color_data = 12'b111111111111;
            11'b00100001101: color_data = 12'b000000000000;
            11'b00100001110: color_data = 12'b000000000000;
            11'b00100001111: color_data = 12'b000000000000;
            11'b00100010000: color_data = 12'b111111111111;
            11'b00100010001: color_data = 12'b111111111111;
            11'b00100010010: color_data = 12'b111111111111;
            11'b00100010011: color_data = 12'b111111111111;
            11'b00100010100: color_data = 12'b111111111111;
            11'b00100010101: color_data = 12'b111111111111;
            11'b00100010110: color_data = 12'b111111111111;
            11'b00100010111: color_data = 12'b111111111111;
            11'b00100011000: color_data = 12'b111111111111;
            11'b00100011001: color_data = 12'b111111111111;
            11'b00100011010: color_data = 12'b111111111111;
            11'b00100011011: color_data = 12'b111111111111;
            11'b00100011100: color_data = 12'b111111111111;
            11'b00100011101: color_data = 12'b111111111111;
            11'b00100011110: color_data = 12'b111111111111;
            11'b00100011111: color_data = 12'b111111111111;
            11'b00100100000: color_data = 12'b111111111111;
            11'b00100100001: color_data = 12'b111111111111;
            11'b00100100010: color_data = 12'b111111111111;
            11'b00100100011: color_data = 12'b111111111111;
            11'b00100100100: color_data = 12'b111111111111;
            11'b00100100101: color_data = 12'b111111111111;
            11'b00100100110: color_data = 12'b111111111111;
            11'b00100100111: color_data = 12'b111111111111;
            11'b00100101000: color_data = 12'b111111111111;
            11'b00100101001: color_data = 12'b111111111111;
            11'b00100101010: color_data = 12'b111111111111;
            11'b00100101011: color_data = 12'b111111111111;
            11'b00100101100: color_data = 12'b000000000000;
            11'b00100101101: color_data = 12'b000000000000;
            11'b00100101110: color_data = 12'b111111111111;
            11'b00100101111: color_data = 12'b111111111111;
            11'b00100110000: color_data = 12'b111111111111;
            11'b00100110001: color_data = 12'b111111111111;
            11'b00100110010: color_data = 12'b111111111111;
            11'b00100110011: color_data = 12'b111111111111;
            11'b00100110100: color_data = 12'b111111111111;
            11'b00100110101: color_data = 12'b111111111111;
            11'b00100110110: color_data = 12'b111111111111;
            11'b00100110111: color_data = 12'b111111111111;
            11'b00100111000: color_data = 12'b111111111111;
            11'b00100111001: color_data = 12'b111111111111;
            11'b00100111010: color_data = 12'b111111111111;
            11'b00100111011: color_data = 12'b111111111111;
            11'b00100111100: color_data = 12'b111111111111;
            11'b00100111101: color_data = 12'b111111111111;
            11'b00100111110: color_data = 12'b111111111111;
            11'b00100111111: color_data = 12'b111111111111;
            11'b00101000000: color_data = 12'b111111111111;
            11'b00101000001: color_data = 12'b111111111111;
            11'b00101000010: color_data = 12'b111111111111;
            11'b00101000011: color_data = 12'b111111111111;
            11'b00101000100: color_data = 12'b111111111111;
            11'b00101000101: color_data = 12'b111111111111;
            11'b00101000110: color_data = 12'b111111111111;
            11'b00101000111: color_data = 12'b111111111111;
            11'b00101001000: color_data = 12'b111111111111;
            11'b00101001001: color_data = 12'b000000000000;
            11'b00101001010: color_data = 12'b000000000000;
            11'b00101001011: color_data = 12'b000000000000;
            11'b00101001100: color_data = 12'b111111111111;
            11'b00101001101: color_data = 12'b111111111111;
            11'b00110000000: color_data = 12'b111111111111;
            11'b00110000001: color_data = 12'b000000000000;
            11'b00110000010: color_data = 12'b000000000000;
            11'b00110000011: color_data = 12'b000000000000;
            11'b00110000100: color_data = 12'b000000000000;
            11'b00110000101: color_data = 12'b111111111111;
            11'b00110000110: color_data = 12'b111111111111;
            11'b00110000111: color_data = 12'b111111111111;
            11'b00110001000: color_data = 12'b111111111111;
            11'b00110001001: color_data = 12'b111111111111;
            11'b00110001010: color_data = 12'b111111111111;
            11'b00110001011: color_data = 12'b111111111111;
            11'b00110001100: color_data = 12'b000000000000;
            11'b00110001101: color_data = 12'b000000000000;
            11'b00110001110: color_data = 12'b111111111111;
            11'b00110001111: color_data = 12'b000000000000;
            11'b00110010000: color_data = 12'b000000000000;
            11'b00110010001: color_data = 12'b111111111111;
            11'b00110010010: color_data = 12'b111111111111;
            11'b00110010011: color_data = 12'b111111111111;
            11'b00110010100: color_data = 12'b111111111111;
            11'b00110010101: color_data = 12'b111111111111;
            11'b00110010110: color_data = 12'b111111111111;
            11'b00110010111: color_data = 12'b111111111111;
            11'b00110011000: color_data = 12'b111111111111;
            11'b00110011001: color_data = 12'b111111111111;
            11'b00110011010: color_data = 12'b111111111111;
            11'b00110011011: color_data = 12'b111111111111;
            11'b00110011100: color_data = 12'b111111111111;
            11'b00110011101: color_data = 12'b111111111111;
            11'b00110011110: color_data = 12'b111111111111;
            11'b00110011111: color_data = 12'b000000000000;
            11'b00110100000: color_data = 12'b000000000000;
            11'b00110100001: color_data = 12'b000000000000;
            11'b00110100010: color_data = 12'b000000000000;
            11'b00110100011: color_data = 12'b111111111111;
            11'b00110100100: color_data = 12'b111111111111;
            11'b00110100101: color_data = 12'b111111111111;
            11'b00110100110: color_data = 12'b111111111111;
            11'b00110100111: color_data = 12'b111111111111;
            11'b00110101000: color_data = 12'b111111111111;
            11'b00110101001: color_data = 12'b111111111111;
            11'b00110101010: color_data = 12'b000000000000;
            11'b00110101011: color_data = 12'b000000000000;
            11'b00110101100: color_data = 12'b000000000000;
            11'b00110101101: color_data = 12'b000000000000;
            11'b00110101110: color_data = 12'b111111111111;
            11'b00110101111: color_data = 12'b111111111111;
            11'b00110110000: color_data = 12'b111111111111;
            11'b00110110001: color_data = 12'b111111111111;
            11'b00110110010: color_data = 12'b111111111111;
            11'b00110110011: color_data = 12'b111111111111;
            11'b00110110100: color_data = 12'b111111111111;
            11'b00110110101: color_data = 12'b111111111111;
            11'b00110110110: color_data = 12'b111111111111;
            11'b00110110111: color_data = 12'b111111111111;
            11'b00110111000: color_data = 12'b111111111111;
            11'b00110111001: color_data = 12'b111111111111;
            11'b00110111010: color_data = 12'b111111111111;
            11'b00110111011: color_data = 12'b111111111111;
            11'b00110111100: color_data = 12'b111111111111;
            11'b00110111101: color_data = 12'b000000000000;
            11'b00110111110: color_data = 12'b000000000000;
            11'b00110111111: color_data = 12'b000000000000;
            11'b00111000000: color_data = 12'b000000000000;
            11'b00111000001: color_data = 12'b111111111111;
            11'b00111000010: color_data = 12'b111111111111;
            11'b00111000011: color_data = 12'b111111111111;
            11'b00111000100: color_data = 12'b111111111111;
            11'b00111000101: color_data = 12'b111111111111;
            11'b00111000110: color_data = 12'b111111111111;
            11'b00111000111: color_data = 12'b111111111111;
            11'b00111001000: color_data = 12'b000000000000;
            11'b00111001001: color_data = 12'b000000000000;
            11'b00111001010: color_data = 12'b111111111111;
            11'b00111001011: color_data = 12'b000000000000;
            11'b00111001100: color_data = 12'b000000000000;
            11'b00111001101: color_data = 12'b111111111111;
            11'b01000000000: color_data = 12'b000000000000;
            11'b01000000001: color_data = 12'b000000000000;
            11'b01000000010: color_data = 12'b111111111111;
            11'b01000000011: color_data = 12'b111111111111;
            11'b01000000100: color_data = 12'b000000000000;
            11'b01000000101: color_data = 12'b000000000000;
            11'b01000000110: color_data = 12'b000000000000;
            11'b01000000111: color_data = 12'b111111111111;
            11'b01000001000: color_data = 12'b000000000000;
            11'b01000001001: color_data = 12'b111111111111;
            11'b01000001010: color_data = 12'b000000000000;
            11'b01000001011: color_data = 12'b000000000000;
            11'b01000001100: color_data = 12'b000000000000;
            11'b01000001101: color_data = 12'b000000000000;
            11'b01000001110: color_data = 12'b111111111111;
            11'b01000001111: color_data = 12'b000000000000;
            11'b01000010000: color_data = 12'b000000000000;
            11'b01000010001: color_data = 12'b111111111111;
            11'b01000010010: color_data = 12'b111111111111;
            11'b01000010011: color_data = 12'b111111111111;
            11'b01000010100: color_data = 12'b111111111111;
            11'b01000010101: color_data = 12'b111111111111;
            11'b01000010110: color_data = 12'b111111111111;
            11'b01000010111: color_data = 12'b111111111111;
            11'b01000011000: color_data = 12'b111111111111;
            11'b01000011001: color_data = 12'b111111111111;
            11'b01000011010: color_data = 12'b111111111111;
            11'b01000011011: color_data = 12'b111111111111;
            11'b01000011100: color_data = 12'b111111111111;
            11'b01000011101: color_data = 12'b111111111111;
            11'b01000011110: color_data = 12'b000000000000;
            11'b01000011111: color_data = 12'b000000000000;
            11'b01000100000: color_data = 12'b111111111111;
            11'b01000100001: color_data = 12'b111111111111;
            11'b01000100010: color_data = 12'b000000000000;
            11'b01000100011: color_data = 12'b000000000000;
            11'b01000100100: color_data = 12'b000000000000;
            11'b01000100101: color_data = 12'b111111111111;
            11'b01000100110: color_data = 12'b000000000000;
            11'b01000100111: color_data = 12'b111111111111;
            11'b01000101000: color_data = 12'b000000000000;
            11'b01000101001: color_data = 12'b000000000000;
            11'b01000101010: color_data = 12'b111111111111;
            11'b01000101011: color_data = 12'b111111111111;
            11'b01000101100: color_data = 12'b000000000000;
            11'b01000101101: color_data = 12'b000000000000;
            11'b01000101110: color_data = 12'b111111111111;
            11'b01000101111: color_data = 12'b111111111111;
            11'b01000110000: color_data = 12'b111111111111;
            11'b01000110001: color_data = 12'b111111111111;
            11'b01000110010: color_data = 12'b111111111111;
            11'b01000110011: color_data = 12'b111111111111;
            11'b01000110100: color_data = 12'b111111111111;
            11'b01000110101: color_data = 12'b111111111111;
            11'b01000110110: color_data = 12'b111111111111;
            11'b01000110111: color_data = 12'b111111111111;
            11'b01000111000: color_data = 12'b111111111111;
            11'b01000111001: color_data = 12'b111111111111;
            11'b01000111010: color_data = 12'b111111111111;
            11'b01000111011: color_data = 12'b111111111111;
            11'b01000111100: color_data = 12'b000000000000;
            11'b01000111101: color_data = 12'b000000000000;
            11'b01000111110: color_data = 12'b111111111111;
            11'b01000111111: color_data = 12'b111111111111;
            11'b01001000000: color_data = 12'b000000000000;
            11'b01001000001: color_data = 12'b000000000000;
            11'b01001000010: color_data = 12'b000000000000;
            11'b01001000011: color_data = 12'b111111111111;
            11'b01001000100: color_data = 12'b000000000000;
            11'b01001000101: color_data = 12'b111111111111;
            11'b01001000110: color_data = 12'b000000000000;
            11'b01001000111: color_data = 12'b000000000000;
            11'b01001001000: color_data = 12'b111111111111;
            11'b01001001001: color_data = 12'b111111111111;
            11'b01001001010: color_data = 12'b111111111111;
            11'b01001001011: color_data = 12'b000000000000;
            11'b01001001100: color_data = 12'b000000000000;
            11'b01001001101: color_data = 12'b111111111111;
            11'b01010000000: color_data = 12'b000000000000;
            11'b01010000001: color_data = 12'b000000000000;
            11'b01010000010: color_data = 12'b000000000000;
            11'b01010000011: color_data = 12'b000000000000;
            11'b01010000100: color_data = 12'b111111111111;
            11'b01010000101: color_data = 12'b111111111111;
            11'b01010000110: color_data = 12'b000000000000;
            11'b01010000111: color_data = 12'b111111111111;
            11'b01010001000: color_data = 12'b000000000000;
            11'b01010001001: color_data = 12'b111111111111;
            11'b01010001010: color_data = 12'b000000000000;
            11'b01010001011: color_data = 12'b111111111111;
            11'b01010001100: color_data = 12'b000000000000;
            11'b01010001101: color_data = 12'b000000000000;
            11'b01010001110: color_data = 12'b111111111111;
            11'b01010001111: color_data = 12'b000000000000;
            11'b01010010000: color_data = 12'b000000000000;
            11'b01010010001: color_data = 12'b111111111111;
            11'b01010010010: color_data = 12'b111111111111;
            11'b01010010011: color_data = 12'b111111111111;
            11'b01010010100: color_data = 12'b111111111111;
            11'b01010010101: color_data = 12'b111111111111;
            11'b01010010110: color_data = 12'b111111111111;
            11'b01010010111: color_data = 12'b111111111111;
            11'b01010011000: color_data = 12'b111111111111;
            11'b01010011001: color_data = 12'b111111111111;
            11'b01010011010: color_data = 12'b111111111111;
            11'b01010011011: color_data = 12'b111111111111;
            11'b01010011100: color_data = 12'b111111111111;
            11'b01010011101: color_data = 12'b111111111111;
            11'b01010011110: color_data = 12'b000000000000;
            11'b01010011111: color_data = 12'b000000000000;
            11'b01010100000: color_data = 12'b000000000000;
            11'b01010100001: color_data = 12'b000000000000;
            11'b01010100010: color_data = 12'b111111111111;
            11'b01010100011: color_data = 12'b111111111111;
            11'b01010100100: color_data = 12'b000000000000;
            11'b01010100101: color_data = 12'b111111111111;
            11'b01010100110: color_data = 12'b000000000000;
            11'b01010100111: color_data = 12'b111111111111;
            11'b01010101000: color_data = 12'b000000000000;
            11'b01010101001: color_data = 12'b111111111111;
            11'b01010101010: color_data = 12'b111111111111;
            11'b01010101011: color_data = 12'b111111111111;
            11'b01010101100: color_data = 12'b000000000000;
            11'b01010101101: color_data = 12'b000000000000;
            11'b01010101110: color_data = 12'b111111111111;
            11'b01010101111: color_data = 12'b111111111111;
            11'b01010110000: color_data = 12'b111111111111;
            11'b01010110001: color_data = 12'b111111111111;
            11'b01010110010: color_data = 12'b111111111111;
            11'b01010110011: color_data = 12'b111111111111;
            11'b01010110100: color_data = 12'b111111111111;
            11'b01010110101: color_data = 12'b111111111111;
            11'b01010110110: color_data = 12'b111111111111;
            11'b01010110111: color_data = 12'b111111111111;
            11'b01010111000: color_data = 12'b111111111111;
            11'b01010111001: color_data = 12'b111111111111;
            11'b01010111010: color_data = 12'b111111111111;
            11'b01010111011: color_data = 12'b111111111111;
            11'b01010111100: color_data = 12'b000000000000;
            11'b01010111101: color_data = 12'b000000000000;
            11'b01010111110: color_data = 12'b000000000000;
            11'b01010111111: color_data = 12'b000000000000;
            11'b01011000000: color_data = 12'b111111111111;
            11'b01011000001: color_data = 12'b111111111111;
            11'b01011000010: color_data = 12'b000000000000;
            11'b01011000011: color_data = 12'b111111111111;
            11'b01011000100: color_data = 12'b000000000000;
            11'b01011000101: color_data = 12'b111111111111;
            11'b01011000110: color_data = 12'b000000000000;
            11'b01011000111: color_data = 12'b111111111111;
            11'b01011001000: color_data = 12'b111111111111;
            11'b01011001001: color_data = 12'b111111111111;
            11'b01011001010: color_data = 12'b000000000000;
            11'b01011001011: color_data = 12'b000000000000;
            11'b01011001100: color_data = 12'b111111111111;
            11'b01011001101: color_data = 12'b111111111111;
            11'b01100000000: color_data = 12'b111111111111;
            11'b01100000001: color_data = 12'b111111111111;
            11'b01100000010: color_data = 12'b000000000000;
            11'b01100000011: color_data = 12'b000000000000;
            11'b01100000100: color_data = 12'b000000000000;
            11'b01100000101: color_data = 12'b111111111111;
            11'b01100000110: color_data = 12'b000000000000;
            11'b01100000111: color_data = 12'b000000000000;
            11'b01100001000: color_data = 12'b000000000000;
            11'b01100001001: color_data = 12'b000000000000;
            11'b01100001010: color_data = 12'b000000000000;
            11'b01100001011: color_data = 12'b111111111111;
            11'b01100001100: color_data = 12'b000000000000;
            11'b01100001101: color_data = 12'b000000000000;
            11'b01100001110: color_data = 12'b111111111111;
            11'b01100001111: color_data = 12'b000000000000;
            11'b01100010000: color_data = 12'b000000000000;
            11'b01100010001: color_data = 12'b111111111111;
            11'b01100010010: color_data = 12'b111111111111;
            11'b01100010011: color_data = 12'b111111111111;
            11'b01100010100: color_data = 12'b111111111111;
            11'b01100010101: color_data = 12'b111111111111;
            11'b01100010110: color_data = 12'b111111111111;
            11'b01100010111: color_data = 12'b111111111111;
            11'b01100011000: color_data = 12'b111111111111;
            11'b01100011001: color_data = 12'b111111111111;
            11'b01100011010: color_data = 12'b111111111111;
            11'b01100011011: color_data = 12'b111111111111;
            11'b01100011100: color_data = 12'b111111111111;
            11'b01100011101: color_data = 12'b111111111111;
            11'b01100011110: color_data = 12'b111111111111;
            11'b01100011111: color_data = 12'b111111111111;
            11'b01100100000: color_data = 12'b000000000000;
            11'b01100100001: color_data = 12'b000000000000;
            11'b01100100010: color_data = 12'b000000000000;
            11'b01100100011: color_data = 12'b111111111111;
            11'b01100100100: color_data = 12'b000000000000;
            11'b01100100101: color_data = 12'b000000000000;
            11'b01100100110: color_data = 12'b000000000000;
            11'b01100100111: color_data = 12'b000000000000;
            11'b01100101000: color_data = 12'b000000000000;
            11'b01100101001: color_data = 12'b111111111111;
            11'b01100101010: color_data = 12'b111111111111;
            11'b01100101011: color_data = 12'b111111111111;
            11'b01100101100: color_data = 12'b000000000000;
            11'b01100101101: color_data = 12'b000000000000;
            11'b01100101110: color_data = 12'b111111111111;
            11'b01100101111: color_data = 12'b111111111111;
            11'b01100110000: color_data = 12'b111111111111;
            11'b01100110001: color_data = 12'b111111111111;
            11'b01100110010: color_data = 12'b111111111111;
            11'b01100110011: color_data = 12'b111111111111;
            11'b01100110100: color_data = 12'b111111111111;
            11'b01100110101: color_data = 12'b111111111111;
            11'b01100110110: color_data = 12'b111111111111;
            11'b01100110111: color_data = 12'b111111111111;
            11'b01100111000: color_data = 12'b111111111111;
            11'b01100111001: color_data = 12'b111111111111;
            11'b01100111010: color_data = 12'b111111111111;
            11'b01100111011: color_data = 12'b111111111111;
            11'b01100111100: color_data = 12'b111111111111;
            11'b01100111101: color_data = 12'b111111111111;
            11'b01100111110: color_data = 12'b000000000000;
            11'b01100111111: color_data = 12'b000000000000;
            11'b01101000000: color_data = 12'b000000000000;
            11'b01101000001: color_data = 12'b111111111111;
            11'b01101000010: color_data = 12'b000000000000;
            11'b01101000011: color_data = 12'b000000000000;
            11'b01101000100: color_data = 12'b000000000000;
            11'b01101000101: color_data = 12'b000000000000;
            11'b01101000110: color_data = 12'b000000000000;
            11'b01101000111: color_data = 12'b111111111111;
            11'b01101001000: color_data = 12'b111111111111;
            11'b01101001001: color_data = 12'b000000000000;
            11'b01101001010: color_data = 12'b000000000000;
            11'b01101001011: color_data = 12'b111111111111;
            11'b01101001100: color_data = 12'b111111111111;
            11'b01101001101: color_data = 12'b111111111111;
            11'b01110000000: color_data = 12'b000000000000;
            11'b01110000001: color_data = 12'b111111111111;
            11'b01110000010: color_data = 12'b111111111111;
            11'b01110000011: color_data = 12'b000000000000;
            11'b01110000100: color_data = 12'b000000000000;
            11'b01110000101: color_data = 12'b111111111111;
            11'b01110000110: color_data = 12'b111111111111;
            11'b01110000111: color_data = 12'b000000000000;
            11'b01110001000: color_data = 12'b000000000000;
            11'b01110001001: color_data = 12'b000000000000;
            11'b01110001010: color_data = 12'b000000000000;
            11'b01110001011: color_data = 12'b111111111111;
            11'b01110001100: color_data = 12'b000000000000;
            11'b01110001101: color_data = 12'b000000000000;
            11'b01110001110: color_data = 12'b111111111111;
            11'b01110001111: color_data = 12'b000000000000;
            11'b01110010000: color_data = 12'b000000000000;
            11'b01110010001: color_data = 12'b111111111111;
            11'b01110010010: color_data = 12'b111111111111;
            11'b01110010011: color_data = 12'b111111111111;
            11'b01110010100: color_data = 12'b111111111111;
            11'b01110010101: color_data = 12'b111111111111;
            11'b01110010110: color_data = 12'b111111111111;
            11'b01110010111: color_data = 12'b111111111111;
            11'b01110011000: color_data = 12'b111111111111;
            11'b01110011001: color_data = 12'b111111111111;
            11'b01110011010: color_data = 12'b111111111111;
            11'b01110011011: color_data = 12'b111111111111;
            11'b01110011100: color_data = 12'b111111111111;
            11'b01110011101: color_data = 12'b111111111111;
            11'b01110011110: color_data = 12'b000000000000;
            11'b01110011111: color_data = 12'b111111111111;
            11'b01110100000: color_data = 12'b111111111111;
            11'b01110100001: color_data = 12'b000000000000;
            11'b01110100010: color_data = 12'b000000000000;
            11'b01110100011: color_data = 12'b111111111111;
            11'b01110100100: color_data = 12'b111111111111;
            11'b01110100101: color_data = 12'b000000000000;
            11'b01110100110: color_data = 12'b000000000000;
            11'b01110100111: color_data = 12'b000000000000;
            11'b01110101000: color_data = 12'b000000000000;
            11'b01110101001: color_data = 12'b111111111111;
            11'b01110101010: color_data = 12'b111111111111;
            11'b01110101011: color_data = 12'b111111111111;
            11'b01110101100: color_data = 12'b000000000000;
            11'b01110101101: color_data = 12'b000000000000;
            11'b01110101110: color_data = 12'b111111111111;
            11'b01110101111: color_data = 12'b111111111111;
            11'b01110110000: color_data = 12'b111111111111;
            11'b01110110001: color_data = 12'b111111111111;
            11'b01110110010: color_data = 12'b111111111111;
            11'b01110110011: color_data = 12'b111111111111;
            11'b01110110100: color_data = 12'b111111111111;
            11'b01110110101: color_data = 12'b111111111111;
            11'b01110110110: color_data = 12'b111111111111;
            11'b01110110111: color_data = 12'b111111111111;
            11'b01110111000: color_data = 12'b111111111111;
            11'b01110111001: color_data = 12'b111111111111;
            11'b01110111010: color_data = 12'b111111111111;
            11'b01110111011: color_data = 12'b111111111111;
            11'b01110111100: color_data = 12'b000000000000;
            11'b01110111101: color_data = 12'b111111111111;
            11'b01110111110: color_data = 12'b111111111111;
            11'b01110111111: color_data = 12'b000000000000;
            11'b01111000000: color_data = 12'b000000000000;
            11'b01111000001: color_data = 12'b111111111111;
            11'b01111000010: color_data = 12'b111111111111;
            11'b01111000011: color_data = 12'b000000000000;
            11'b01111000100: color_data = 12'b000000000000;
            11'b01111000101: color_data = 12'b000000000000;
            11'b01111000110: color_data = 12'b000000000000;
            11'b01111000111: color_data = 12'b111111111111;
            11'b01111001000: color_data = 12'b000000000000;
            11'b01111001001: color_data = 12'b000000000000;
            11'b01111001010: color_data = 12'b111111111111;
            11'b01111001011: color_data = 12'b000000000000;
            11'b01111001100: color_data = 12'b000000000000;
            11'b01111001101: color_data = 12'b111111111111;
            11'b10000000000: color_data = 12'b000000000000;
            11'b10000000001: color_data = 12'b000000000000;
            11'b10000000010: color_data = 12'b000000000000;
            11'b10000000011: color_data = 12'b000000000000;
            11'b10000000100: color_data = 12'b111111111111;
            11'b10000000101: color_data = 12'b111111111111;
            11'b10000000110: color_data = 12'b111111111111;
            11'b10000000111: color_data = 12'b000000000000;
            11'b10000001000: color_data = 12'b111111111111;
            11'b10000001001: color_data = 12'b000000000000;
            11'b10000001010: color_data = 12'b111111111111;
            11'b10000001011: color_data = 12'b111111111111;
            11'b10000001100: color_data = 12'b111111111111;
            11'b10000001101: color_data = 12'b000000000000;
            11'b10000001110: color_data = 12'b000000000000;
            11'b10000001111: color_data = 12'b000000000000;
            11'b10000010000: color_data = 12'b111111111111;
            11'b10000010001: color_data = 12'b111111111111;
            11'b10000010010: color_data = 12'b111111111111;
            11'b10000010011: color_data = 12'b111111111111;
            11'b10000010100: color_data = 12'b000000000000;
            11'b10000010101: color_data = 12'b000000000000;
            11'b10000010110: color_data = 12'b111111111111;
            11'b10000010111: color_data = 12'b111111111111;
            11'b10000011000: color_data = 12'b111111111111;
            11'b10000011001: color_data = 12'b111111111111;
            11'b10000011010: color_data = 12'b111111111111;
            11'b10000011011: color_data = 12'b111111111111;
            11'b10000011100: color_data = 12'b111111111111;
            11'b10000011101: color_data = 12'b111111111111;
            11'b10000011110: color_data = 12'b000000000000;
            11'b10000011111: color_data = 12'b000000000000;
            11'b10000100000: color_data = 12'b000000000000;
            11'b10000100001: color_data = 12'b000000000000;
            11'b10000100010: color_data = 12'b111111111111;
            11'b10000100011: color_data = 12'b111111111111;
            11'b10000100100: color_data = 12'b111111111111;
            11'b10000100101: color_data = 12'b000000000000;
            11'b10000100110: color_data = 12'b111111111111;
            11'b10000100111: color_data = 12'b000000000000;
            11'b10000101000: color_data = 12'b111111111111;
            11'b10000101001: color_data = 12'b111111111111;
            11'b10000101010: color_data = 12'b000000000000;
            11'b10000101011: color_data = 12'b000000000000;
            11'b10000101100: color_data = 12'b000000000000;
            11'b10000101101: color_data = 12'b000000000000;
            11'b10000101110: color_data = 12'b000000000000;
            11'b10000101111: color_data = 12'b000000000000;
            11'b10000110000: color_data = 12'b111111111111;
            11'b10000110001: color_data = 12'b111111111111;
            11'b10000110010: color_data = 12'b000000000000;
            11'b10000110011: color_data = 12'b000000000000;
            11'b10000110100: color_data = 12'b111111111111;
            11'b10000110101: color_data = 12'b111111111111;
            11'b10000110110: color_data = 12'b111111111111;
            11'b10000110111: color_data = 12'b111111111111;
            11'b10000111000: color_data = 12'b111111111111;
            11'b10000111001: color_data = 12'b111111111111;
            11'b10000111010: color_data = 12'b111111111111;
            11'b10000111011: color_data = 12'b111111111111;
            11'b10000111100: color_data = 12'b000000000000;
            11'b10000111101: color_data = 12'b000000000000;
            11'b10000111110: color_data = 12'b000000000000;
            11'b10000111111: color_data = 12'b000000000000;
            11'b10001000000: color_data = 12'b111111111111;
            11'b10001000001: color_data = 12'b111111111111;
            11'b10001000010: color_data = 12'b111111111111;
            11'b10001000011: color_data = 12'b000000000000;
            11'b10001000100: color_data = 12'b111111111111;
            11'b10001000101: color_data = 12'b000000000000;
            11'b10001000110: color_data = 12'b111111111111;
            11'b10001000111: color_data = 12'b111111111111;
            11'b10001001000: color_data = 12'b000000000000;
            11'b10001001001: color_data = 12'b000000000000;
            11'b10001001010: color_data = 12'b000000000000;
            11'b10001001011: color_data = 12'b000000000000;
            11'b10001001100: color_data = 12'b000000000000;
            11'b10001001101: color_data = 12'b111111111111;
            11'b10010000000: color_data = 12'b111111111111;
            11'b10010000001: color_data = 12'b111111111111;
            11'b10010000010: color_data = 12'b111111111111;
            11'b10010000011: color_data = 12'b111111111111;
            11'b10010000100: color_data = 12'b111111111111;
            11'b10010000101: color_data = 12'b111111111111;
            11'b10010000110: color_data = 12'b111111111111;
            11'b10010000111: color_data = 12'b111111111111;
            11'b10010001000: color_data = 12'b111111111111;
            11'b10010001001: color_data = 12'b111111111111;
            11'b10010001010: color_data = 12'b111111111111;
            11'b10010001011: color_data = 12'b111111111111;
            11'b10010001100: color_data = 12'b111111111111;
            11'b10010001101: color_data = 12'b111111111111;
            11'b10010001110: color_data = 12'b111111111111;
            11'b10010001111: color_data = 12'b111111111111;
            11'b10010010000: color_data = 12'b111111111111;
            11'b10010010001: color_data = 12'b111111111111;
            11'b10010010010: color_data = 12'b111111111111;
            11'b10010010011: color_data = 12'b111111111111;
            11'b10010010100: color_data = 12'b000000000000;
            11'b10010010101: color_data = 12'b111111111111;
            11'b10010010110: color_data = 12'b111111111111;
            11'b10010010111: color_data = 12'b111111111111;
            11'b10010011000: color_data = 12'b111111111111;
            11'b10010011001: color_data = 12'b111111111111;
            11'b10010011010: color_data = 12'b111111111111;
            11'b10010011011: color_data = 12'b111111111111;
            11'b10010011100: color_data = 12'b111111111111;
            11'b10010011101: color_data = 12'b111111111111;
            11'b10010011110: color_data = 12'b111111111111;
            11'b10010011111: color_data = 12'b111111111111;
            11'b10010100000: color_data = 12'b111111111111;
            11'b10010100001: color_data = 12'b111111111111;
            11'b10010100010: color_data = 12'b111111111111;
            11'b10010100011: color_data = 12'b111111111111;
            11'b10010100100: color_data = 12'b111111111111;
            11'b10010100101: color_data = 12'b111111111111;
            11'b10010100110: color_data = 12'b111111111111;
            11'b10010100111: color_data = 12'b111111111111;
            11'b10010101000: color_data = 12'b111111111111;
            11'b10010101001: color_data = 12'b111111111111;
            11'b10010101010: color_data = 12'b111111111111;
            11'b10010101011: color_data = 12'b111111111111;
            11'b10010101100: color_data = 12'b111111111111;
            11'b10010101101: color_data = 12'b111111111111;
            11'b10010101110: color_data = 12'b111111111111;
            11'b10010101111: color_data = 12'b111111111111;
            11'b10010110000: color_data = 12'b111111111111;
            11'b10010110001: color_data = 12'b111111111111;
            11'b10010110010: color_data = 12'b000000000000;
            11'b10010110011: color_data = 12'b111111111111;
            11'b10010110100: color_data = 12'b111111111111;
            11'b10010110101: color_data = 12'b111111111111;
            11'b10010110110: color_data = 12'b111111111111;
            11'b10010110111: color_data = 12'b111111111111;
            11'b10010111000: color_data = 12'b111111111111;
            11'b10010111001: color_data = 12'b111111111111;
            11'b10010111010: color_data = 12'b111111111111;
            11'b10010111011: color_data = 12'b111111111111;
            11'b10010111100: color_data = 12'b111111111111;
            11'b10010111101: color_data = 12'b111111111111;
            11'b10010111110: color_data = 12'b111111111111;
            11'b10010111111: color_data = 12'b111111111111;
            11'b10011000000: color_data = 12'b111111111111;
            11'b10011000001: color_data = 12'b111111111111;
            11'b10011000010: color_data = 12'b111111111111;
            11'b10011000011: color_data = 12'b111111111111;
            11'b10011000100: color_data = 12'b111111111111;
            11'b10011000101: color_data = 12'b111111111111;
            11'b10011000110: color_data = 12'b111111111111;
            11'b10011000111: color_data = 12'b111111111111;
            11'b10011001000: color_data = 12'b111111111111;
            11'b10011001001: color_data = 12'b111111111111;
            11'b10011001010: color_data = 12'b111111111111;
            11'b10011001011: color_data = 12'b111111111111;
            11'b10011001100: color_data = 12'b111111111111;
            11'b10011001101: color_data = 12'b111111111111;
            11'b10100000000: color_data = 12'b111111111111;
            11'b10100000001: color_data = 12'b111111111111;
            11'b10100000010: color_data = 12'b111111111111;
            11'b10100000011: color_data = 12'b111111111111;
            11'b10100000100: color_data = 12'b111111111111;
            11'b10100000101: color_data = 12'b111111111111;
            11'b10100000110: color_data = 12'b111111111111;
            11'b10100000111: color_data = 12'b111111111111;
            11'b10100001000: color_data = 12'b111111111111;
            11'b10100001001: color_data = 12'b111111111111;
            11'b10100001010: color_data = 12'b111111111111;
            11'b10100001011: color_data = 12'b111111111111;
            11'b10100001100: color_data = 12'b111111111111;
            11'b10100001101: color_data = 12'b111111111111;
            11'b10100001110: color_data = 12'b111111111111;
            11'b10100001111: color_data = 12'b111111111111;
            11'b10100010000: color_data = 12'b111111111111;
            11'b10100010001: color_data = 12'b111111111111;
            11'b10100010010: color_data = 12'b111111111111;
            11'b10100010011: color_data = 12'b000000000000;
            11'b10100010100: color_data = 12'b111111111111;
            11'b10100010101: color_data = 12'b111111111111;
            11'b10100010110: color_data = 12'b111111111111;
            11'b10100010111: color_data = 12'b111111111111;
            11'b10100011000: color_data = 12'b111111111111;
            11'b10100011001: color_data = 12'b111111111111;
            11'b10100011010: color_data = 12'b111111111111;
            11'b10100011011: color_data = 12'b111111111111;
            11'b10100011100: color_data = 12'b111111111111;
            11'b10100011101: color_data = 12'b111111111111;
            11'b10100011110: color_data = 12'b111111111111;
            11'b10100011111: color_data = 12'b111111111111;
            11'b10100100000: color_data = 12'b111111111111;
            11'b10100100001: color_data = 12'b111111111111;
            11'b10100100010: color_data = 12'b111111111111;
            11'b10100100011: color_data = 12'b111111111111;
            11'b10100100100: color_data = 12'b111111111111;
            11'b10100100101: color_data = 12'b111111111111;
            11'b10100100110: color_data = 12'b111111111111;
            11'b10100100111: color_data = 12'b111111111111;
            11'b10100101000: color_data = 12'b111111111111;
            11'b10100101001: color_data = 12'b111111111111;
            11'b10100101010: color_data = 12'b111111111111;
            11'b10100101011: color_data = 12'b111111111111;
            11'b10100101100: color_data = 12'b111111111111;
            11'b10100101101: color_data = 12'b111111111111;
            11'b10100101110: color_data = 12'b111111111111;
            11'b10100101111: color_data = 12'b111111111111;
            11'b10100110000: color_data = 12'b111111111111;
            11'b10100110001: color_data = 12'b000000000000;
            11'b10100110010: color_data = 12'b111111111111;
            11'b10100110011: color_data = 12'b111111111111;
            11'b10100110100: color_data = 12'b111111111111;
            11'b10100110101: color_data = 12'b111111111111;
            11'b10100110110: color_data = 12'b111111111111;
            11'b10100110111: color_data = 12'b111111111111;
            11'b10100111000: color_data = 12'b111111111111;
            11'b10100111001: color_data = 12'b111111111111;
            11'b10100111010: color_data = 12'b111111111111;
            11'b10100111011: color_data = 12'b111111111111;
            11'b10100111100: color_data = 12'b111111111111;
            11'b10100111101: color_data = 12'b111111111111;
            11'b10100111110: color_data = 12'b111111111111;
            11'b10100111111: color_data = 12'b111111111111;
            11'b10101000000: color_data = 12'b111111111111;
            11'b10101000001: color_data = 12'b111111111111;
            11'b10101000010: color_data = 12'b111111111111;
            11'b10101000011: color_data = 12'b111111111111;
            11'b10101000100: color_data = 12'b111111111111;
            11'b10101000101: color_data = 12'b111111111111;
            11'b10101000110: color_data = 12'b111111111111;
            11'b10101000111: color_data = 12'b111111111111;
            11'b10101001000: color_data = 12'b111111111111;
            11'b10101001001: color_data = 12'b111111111111;
            11'b10101001010: color_data = 12'b111111111111;
            11'b10101001011: color_data = 12'b111111111111;
            11'b10101001100: color_data = 12'b111111111111;
            11'b10101001101: color_data = 12'b111111111111;
            default:       color_data = 12'b000000000000;
        endcase
    end
endmodule
