module italian_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=12'b000000000000) && ({row_reg, col_reg}<12'b000000001111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000000001111) && ({row_reg, col_reg}<12'b000000010010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000000010010) && ({row_reg, col_reg}<12'b000000011010)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000000011010) && ({row_reg, col_reg}<12'b000000011110)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000000011110) && ({row_reg, col_reg}<12'b000000100000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000000100000)) color_data = 12'b111100010110;

		if(({row_reg, col_reg}>=12'b000000100001) && ({row_reg, col_reg}<12'b000001010000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000001010000) && ({row_reg, col_reg}<12'b000001010010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000001010010) && ({row_reg, col_reg}<12'b000001011010)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000001011010) && ({row_reg, col_reg}<12'b000001011101)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b000001011101) && ({row_reg, col_reg}<12'b000010000000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000010000000) && ({row_reg, col_reg}<12'b000010000010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000010000010) && ({row_reg, col_reg}<12'b000010000111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000010000111)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b000010001000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000010001001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000010001010) && ({row_reg, col_reg}<12'b000010001110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000010001110) && ({row_reg, col_reg}<12'b000010010001)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b000010010001) && ({row_reg, col_reg}<12'b000011000000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000011000000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000011000001) && ({row_reg, col_reg}<12'b000011000111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000011000111)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b000011001000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000011001001) && ({row_reg, col_reg}<12'b000011001101)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000011001101) && ({row_reg, col_reg}<12'b000011011110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000011011110) && ({row_reg, col_reg}<12'b000011100011)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b000011100011) && ({row_reg, col_reg}<12'b000100000110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000100000110) && ({row_reg, col_reg}<12'b000100001101)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000100001101) && ({row_reg, col_reg}<12'b000100010000)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}>=12'b000100010000) && ({row_reg, col_reg}<12'b000100010010)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000100010010) && ({row_reg, col_reg}<12'b000100010100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000100010100) && ({row_reg, col_reg}<12'b000100011011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000100011011)) color_data = 12'b111100010110;
		if(({row_reg, col_reg}>=12'b000100011100) && ({row_reg, col_reg}<12'b000100011110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000100011110) && ({row_reg, col_reg}<12'b000100100011)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b000100100011) && ({row_reg, col_reg}<12'b000101000110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000101000110) && ({row_reg, col_reg}<12'b000101001001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000101001001) && ({row_reg, col_reg}<12'b000101001100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000101001100) && ({row_reg, col_reg}<12'b000101010000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000101010000) && ({row_reg, col_reg}<12'b000101010010)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000101010010) && ({row_reg, col_reg}<12'b000101010100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000101010100) && ({row_reg, col_reg}<12'b000101011000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000101011000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000101011001) && ({row_reg, col_reg}<12'b000101011011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000101011011)) color_data = 12'b111100010110;
		if(({row_reg, col_reg}>=12'b000101011100) && ({row_reg, col_reg}<12'b000101011111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000101011111) && ({row_reg, col_reg}<12'b000101100011)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b000101100011) && ({row_reg, col_reg}<12'b000110000010)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000110000010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000110000011) && ({row_reg, col_reg}<12'b000110001100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000110001100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000110001101) && ({row_reg, col_reg}<12'b000110010001)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b000110010001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000110010010) && ({row_reg, col_reg}<12'b000110010111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000110010111) && ({row_reg, col_reg}<12'b000110011010)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b000110011010) && ({row_reg, col_reg}<12'b000111000001)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000111000001) && ({row_reg, col_reg}<12'b000111000011)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000111000011) && ({row_reg, col_reg}<12'b000111001011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b000111001011)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b000111001100)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b000111001101)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b000111001110)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==12'b000111001111)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==12'b000111010000)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b000111010001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b000111010010) && ({row_reg, col_reg}<12'b000111010111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b000111010111) && ({row_reg, col_reg}<12'b000111011011)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b000111011011) && ({row_reg, col_reg}<12'b001000000101)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001000000101)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001000000110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001000000111)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001000001000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001000001001)) color_data = 12'b111100010110;
		if(({row_reg, col_reg}==12'b001000001010)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001000001011)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001000001100)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b001000001101)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==12'b001000001110)) color_data = 12'b011100110101;
		if(({row_reg, col_reg}==12'b001000001111)) color_data = 12'b100000100100;
		if(({row_reg, col_reg}==12'b001000010000)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}>=12'b001000010001) && ({row_reg, col_reg}<12'b001000010111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b001000010111) && ({row_reg, col_reg}<12'b001000011010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001000011010) && ({row_reg, col_reg}<12'b001000100000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b001000100000) && ({row_reg, col_reg}<12'b001000100010)) color_data = 12'b111100010110;
		if(({row_reg, col_reg}>=12'b001000100010) && ({row_reg, col_reg}<12'b001000100100)) color_data = 12'b111000010110;

		if(({row_reg, col_reg}==12'b001000100100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001001000000) && ({row_reg, col_reg}<12'b001001000101)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b001001000101) && ({row_reg, col_reg}<12'b001001001011)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b001001001011)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b001001001100)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==12'b001001001101)) color_data = 12'b100000110101;
		if(({row_reg, col_reg}==12'b001001001110)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==12'b001001001111)) color_data = 12'b011100110101;
		if(({row_reg, col_reg}==12'b001001010000)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b001001010001)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001001010010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001001010011) && ({row_reg, col_reg}<12'b001001100000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b001001100000) && ({row_reg, col_reg}<12'b001001100011)) color_data = 12'b111100010110;

		if(({row_reg, col_reg}>=12'b001001100011) && ({row_reg, col_reg}<12'b001010000000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001010000000)) color_data = 12'b111100010110;
		if(({row_reg, col_reg}>=12'b001010000001) && ({row_reg, col_reg}<12'b001010000011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001010000011)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001010000100)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b001010000101)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==12'b001010000110)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==12'b001010000111)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}>=12'b001010001000) && ({row_reg, col_reg}<12'b001010001010)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==12'b001010001010)) color_data = 12'b100101000110;
		if(({row_reg, col_reg}==12'b001010001011)) color_data = 12'b100001000110;
		if(({row_reg, col_reg}>=12'b001010001100) && ({row_reg, col_reg}<12'b001010001110)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==12'b001010001110)) color_data = 12'b011001010110;
		if(({row_reg, col_reg}==12'b001010001111)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}==12'b001010010000)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}>=12'b001010010001) && ({row_reg, col_reg}<12'b001010010011)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001010010011) && ({row_reg, col_reg}<12'b001010011110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b001010011110) && ({row_reg, col_reg}<12'b001010100000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001010100000)) color_data = 12'b111100010110;
		if(({row_reg, col_reg}>=12'b001010100001) && ({row_reg, col_reg}<12'b001010100100)) color_data = 12'b111000010110;

		if(({row_reg, col_reg}==12'b001010100100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001011000000)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}==12'b001011000001)) color_data = 12'b110100010110;
		if(({row_reg, col_reg}==12'b001011000010)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b001011000011)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==12'b001011000100)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==12'b001011000101)) color_data = 12'b101001010110;
		if(({row_reg, col_reg}>=12'b001011000110) && ({row_reg, col_reg}<12'b001011001001)) color_data = 12'b100101010110;
		if(({row_reg, col_reg}==12'b001011001001)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==12'b001011001010)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==12'b001011001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b001011001100)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==12'b001011001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001011001110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==12'b001011001111)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==12'b001011010000)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==12'b001011010001)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b001011010010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001011010011) && ({row_reg, col_reg}<12'b001011011110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b001011011110) && ({row_reg, col_reg}<12'b001011100001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001011100001) && ({row_reg, col_reg}<12'b001011100011)) color_data = 12'b111000010110;

		if(({row_reg, col_reg}>=12'b001011100011) && ({row_reg, col_reg}<12'b001100000000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001100000000)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b001100000001)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b001100000010)) color_data = 12'b101101010111;
		if(({row_reg, col_reg}==12'b001100000011)) color_data = 12'b101001111000;
		if(({row_reg, col_reg}==12'b001100000100)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==12'b001100000101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b001100000110)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=12'b001100000111) && ({row_reg, col_reg}<12'b001100001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=12'b001100001011) && ({row_reg, col_reg}<12'b001100001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001100001111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==12'b001100010000)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==12'b001100010001)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==12'b001100010010)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}>=12'b001100010011) && ({row_reg, col_reg}<12'b001100010110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b001100010110) && ({row_reg, col_reg}<12'b001100011000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001100011000) && ({row_reg, col_reg}<12'b001100011010)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b001100011010) && ({row_reg, col_reg}<12'b001100011100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001100011100) && ({row_reg, col_reg}<12'b001100011110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b001100011110) && ({row_reg, col_reg}<12'b001100100000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001100100000) && ({row_reg, col_reg}<12'b001100100010)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}>=12'b001100100010) && ({row_reg, col_reg}<12'b001100100100)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}==12'b001100100100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001101000000)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b001101000001)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}==12'b001101000010)) color_data = 12'b101101101000;
		if(({row_reg, col_reg}==12'b001101000011)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==12'b001101000100)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==12'b001101000101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b001101000110) && ({row_reg, col_reg}<12'b001101001000)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b001101001000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=12'b001101001001) && ({row_reg, col_reg}<12'b001101001011)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}>=12'b001101001011) && ({row_reg, col_reg}<12'b001101010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001101010000)) color_data = 12'b011001010110;
		if(({row_reg, col_reg}==12'b001101010001)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==12'b001101010010)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==12'b001101010011)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b001101010100)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}>=12'b001101010101) && ({row_reg, col_reg}<12'b001101011000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001101011000) && ({row_reg, col_reg}<12'b001101011010)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001101011010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001101011011) && ({row_reg, col_reg}<12'b001101011110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001101011110)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001101011111) && ({row_reg, col_reg}<12'b001101100100)) color_data = 12'b110100100110;

		if(({row_reg, col_reg}>=12'b001101100100) && ({row_reg, col_reg}<12'b001110000001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001110000001)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b001110000010)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==12'b001110000011)) color_data = 12'b110001111000;
		if(({row_reg, col_reg}==12'b001110000100)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==12'b001110000101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b001110000110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b001110000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001110001000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b001110001001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b001110001010)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}>=12'b001110001011) && ({row_reg, col_reg}<12'b001110001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001110001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001110001110)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==12'b001110001111)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==12'b001110010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001110010001)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==12'b001110010010)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}==12'b001110010011)) color_data = 12'b100101000101;
		if(({row_reg, col_reg}==12'b001110010100)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b001110010101)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b001110010110)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001110010111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b001110011000) && ({row_reg, col_reg}<12'b001110011010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b001110011010) && ({row_reg, col_reg}<12'b001110011110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001110011110)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001110011111)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b001110100000)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}>=12'b001110100001) && ({row_reg, col_reg}<12'b001110100011)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b001110100011)) color_data = 12'b110100100110;

		if(({row_reg, col_reg}==12'b001110100100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001111000000)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b001111000001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001111000010)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b001111000011)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==12'b001111000100)) color_data = 12'b101101010111;
		if(({row_reg, col_reg}==12'b001111000101)) color_data = 12'b101001100111;
		if(({row_reg, col_reg}>=12'b001111000110) && ({row_reg, col_reg}<12'b001111001000)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==12'b001111001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b001111001001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==12'b001111001010)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==12'b001111001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b001111001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001111001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001111001110)) color_data = 12'b010101100101;
		if(({row_reg, col_reg}>=12'b001111001111) && ({row_reg, col_reg}<12'b001111010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001111010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001111010011)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==12'b001111010100)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==12'b001111010101)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}>=12'b001111010110) && ({row_reg, col_reg}<12'b001111011001)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b001111011001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001111011010)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001111011011)) color_data = 12'b111100010110;
		if(({row_reg, col_reg}==12'b001111011100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b001111011101)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b001111011110)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b001111011111)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b001111100000)) color_data = 12'b101100010100;
		if(({row_reg, col_reg}==12'b001111100001)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==12'b001111100010)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b001111100011)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}==12'b001111100100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b010000000000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b010000000001) && ({row_reg, col_reg}<12'b010000000011)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}==12'b010000000011)) color_data = 12'b110100100101;
		if(({row_reg, col_reg}==12'b010000000100)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b010000000101)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010000000110)) color_data = 12'b110001010111;
		if(({row_reg, col_reg}==12'b010000000111)) color_data = 12'b110001111000;
		if(({row_reg, col_reg}==12'b010000001000)) color_data = 12'b110010001001;
		if(({row_reg, col_reg}==12'b010000001001)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==12'b010000001010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b010000001011)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==12'b010000001100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b010000001101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==12'b010000001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010000001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010000010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010000010001)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==12'b010000010010)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==12'b010000010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010000010100)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==12'b010000010101)) color_data = 12'b100101000110;
		if(({row_reg, col_reg}==12'b010000010110)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}>=12'b010000010111) && ({row_reg, col_reg}<12'b010000011001)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010000011001)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b010000011010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b010000011011) && ({row_reg, col_reg}<12'b010000011101)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b010000011101)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010000011110)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==12'b010000011111)) color_data = 12'b100000100100;
		if(({row_reg, col_reg}==12'b010000100000)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b010000100001)) color_data = 12'b110100010101;
		if(({row_reg, col_reg}>=12'b010000100010) && ({row_reg, col_reg}<12'b010000100100)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}==12'b010000100100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b010001000000)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b010001000001)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b010001000010)) color_data = 12'b111100010110;
		if(({row_reg, col_reg}>=12'b010001000011) && ({row_reg, col_reg}<12'b010001000101)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b010001000101)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010001000110)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b010001000111)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==12'b010001001000)) color_data = 12'b101001010110;
		if(({row_reg, col_reg}==12'b010001001001)) color_data = 12'b101001100111;
		if(({row_reg, col_reg}==12'b010001001010)) color_data = 12'b100101100110;
		if(({row_reg, col_reg}>=12'b010001001011) && ({row_reg, col_reg}<12'b010001001101)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==12'b010001001101)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==12'b010001001110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==12'b010001001111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==12'b010001010000)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==12'b010001010001)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==12'b010001010010)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==12'b010001010011)) color_data = 12'b001101000011;
		if(({row_reg, col_reg}==12'b010001010100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010001010101)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==12'b010001010110)) color_data = 12'b100001000101;
		if(({row_reg, col_reg}==12'b010001010111)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==12'b010001011000)) color_data = 12'b101000110110;
		if(({row_reg, col_reg}==12'b010001011001)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==12'b010001011010)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==12'b010001011011)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010001011100)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b010001011101)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==12'b010001011110)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}==12'b010001011111)) color_data = 12'b100000100100;
		if(({row_reg, col_reg}==12'b010001100000)) color_data = 12'b110100100101;

		if(({row_reg, col_reg}>=12'b010001100001) && ({row_reg, col_reg}<12'b010010000000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b010010000000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b010010000001) && ({row_reg, col_reg}<12'b010010000011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b010010000011) && ({row_reg, col_reg}<12'b010010000101)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b010010000101)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b010010000110)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010010000111)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b010010001000)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}>=12'b010010001001) && ({row_reg, col_reg}<12'b010010001011)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==12'b010010001011)) color_data = 12'b101001000101;
		if(({row_reg, col_reg}==12'b010010001100)) color_data = 12'b101101010110;
		if(({row_reg, col_reg}==12'b010010001101)) color_data = 12'b101101010111;
		if(({row_reg, col_reg}==12'b010010001110)) color_data = 12'b100001000101;
		if(({row_reg, col_reg}==12'b010010001111)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==12'b010010010000)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}>=12'b010010010001) && ({row_reg, col_reg}<12'b010010010011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==12'b010010010011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010010010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010010010101)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}>=12'b010010010110) && ({row_reg, col_reg}<12'b010010011000)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==12'b010010011000)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==12'b010010011001)) color_data = 12'b100001000101;
		if(({row_reg, col_reg}==12'b010010011010)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==12'b010010011011)) color_data = 12'b101001000101;
		if(({row_reg, col_reg}==12'b010010011100)) color_data = 12'b101001010110;
		if(({row_reg, col_reg}==12'b010010011101)) color_data = 12'b011100110100;
		if(({row_reg, col_reg}==12'b010010011110)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==12'b010010011111)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==12'b010010100000)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010010100001)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b010010100010) && ({row_reg, col_reg}<12'b010011000101)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b010011000101) && ({row_reg, col_reg}<12'b010011000111)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b010011000111)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010011001000)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010011001001)) color_data = 12'b011100000010;
		if(({row_reg, col_reg}==12'b010011001010)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==12'b010011001011)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010011001100)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b010011001101)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==12'b010011001110)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==12'b010011001111)) color_data = 12'b100101010110;
		if(({row_reg, col_reg}>=12'b010011010000) && ({row_reg, col_reg}<12'b010011010010)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==12'b010011010010)) color_data = 12'b100101010110;
		if(({row_reg, col_reg}==12'b010011010011)) color_data = 12'b101001100110;
		if(({row_reg, col_reg}==12'b010011010100)) color_data = 12'b100101010110;
		if(({row_reg, col_reg}==12'b010011010101)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}>=12'b010011010110) && ({row_reg, col_reg}<12'b010011011000)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==12'b010011011000)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}==12'b010011011001)) color_data = 12'b100001000101;
		if(({row_reg, col_reg}==12'b010011011010)) color_data = 12'b101001000101;
		if(({row_reg, col_reg}==12'b010011011011)) color_data = 12'b100101000101;
		if(({row_reg, col_reg}==12'b010011011100)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==12'b010011011101)) color_data = 12'b011000100011;
		if(({row_reg, col_reg}==12'b010011011110)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==12'b010011011111)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b010011100000)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b010011100001) && ({row_reg, col_reg}<12'b010100000011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b010100000011) && ({row_reg, col_reg}<12'b010100000101)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b010100000101)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b010100000110)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b010100000111)) color_data = 12'b110100100101;
		if(({row_reg, col_reg}==12'b010100001000)) color_data = 12'b101000110101;
		if(({row_reg, col_reg}==12'b010100001001)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==12'b010100001010)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b010100001011)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010100001100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b010100001101)) color_data = 12'b110100100101;
		if(({row_reg, col_reg}==12'b010100001110)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b010100001111)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==12'b010100010000)) color_data = 12'b100101000110;
		if(({row_reg, col_reg}==12'b010100010001)) color_data = 12'b100000110101;
		if(({row_reg, col_reg}==12'b010100010010)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==12'b010100010011)) color_data = 12'b110100110101;
		if(({row_reg, col_reg}==12'b010100010100)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b010100010101)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}==12'b010100010110)) color_data = 12'b011100110101;
		if(({row_reg, col_reg}==12'b010100010111)) color_data = 12'b100001000110;
		if(({row_reg, col_reg}==12'b010100011000)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==12'b010100011001)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==12'b010100011010)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b010100011011)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}==12'b010100011100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==12'b010100011101)) color_data = 12'b011100100100;
		if(({row_reg, col_reg}==12'b010100011110)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010100011111)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b010100100000) && ({row_reg, col_reg}<12'b010101000011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b010101000011) && ({row_reg, col_reg}<12'b010101000101)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b010101000101)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010101000110)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b010101000111)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==12'b010101001000)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==12'b010101001001)) color_data = 12'b011000100100;
		if(({row_reg, col_reg}==12'b010101001010)) color_data = 12'b101100100110;
		if(({row_reg, col_reg}==12'b010101001011)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010101001100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b010101001101)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}==12'b010101001110)) color_data = 12'b110100100101;
		if(({row_reg, col_reg}==12'b010101001111)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010101010000)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==12'b010101010001)) color_data = 12'b101000110101;
		if(({row_reg, col_reg}==12'b010101010010)) color_data = 12'b110100100101;
		if(({row_reg, col_reg}==12'b010101010011)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b010101010100)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010101010101)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==12'b010101010110)) color_data = 12'b011100110110;
		if(({row_reg, col_reg}==12'b010101010111)) color_data = 12'b010100100101;
		if(({row_reg, col_reg}==12'b010101011000)) color_data = 12'b101000110110;
		if(({row_reg, col_reg}==12'b010101011001)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010101011010)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010101011011)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010101011100)) color_data = 12'b100000100101;
		if(({row_reg, col_reg}==12'b010101011101)) color_data = 12'b100000100100;
		if(({row_reg, col_reg}==12'b010101011110)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010101011111)) color_data = 12'b111000010101;

		if(({row_reg, col_reg}>=12'b010101100000) && ({row_reg, col_reg}<12'b010110000011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b010110000011)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b010110000100)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010110000101)) color_data = 12'b101100110111;
		if(({row_reg, col_reg}==12'b010110000110)) color_data = 12'b100001001000;
		if(({row_reg, col_reg}==12'b010110000111)) color_data = 12'b011001011000;
		if(({row_reg, col_reg}==12'b010110001000)) color_data = 12'b001101010111;
		if(({row_reg, col_reg}==12'b010110001001)) color_data = 12'b010001000110;
		if(({row_reg, col_reg}==12'b010110001010)) color_data = 12'b100000100110;
		if(({row_reg, col_reg}==12'b010110001011)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010110001100)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}>=12'b010110001101) && ({row_reg, col_reg}<12'b010110001111)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b010110001111)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}>=12'b010110010000) && ({row_reg, col_reg}<12'b010110010010)) color_data = 12'b101000110101;
		if(({row_reg, col_reg}==12'b010110010010)) color_data = 12'b110100100101;
		if(({row_reg, col_reg}==12'b010110010011)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}==12'b010110010100)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b010110010101)) color_data = 12'b100101000111;
		if(({row_reg, col_reg}==12'b010110010110)) color_data = 12'b010001011000;
		if(({row_reg, col_reg}==12'b010110010111)) color_data = 12'b001101000111;
		if(({row_reg, col_reg}==12'b010110011000)) color_data = 12'b011100110111;
		if(({row_reg, col_reg}==12'b010110011001)) color_data = 12'b101100110111;
		if(({row_reg, col_reg}>=12'b010110011010) && ({row_reg, col_reg}<12'b010110011100)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010110011100)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010110011101)) color_data = 12'b100100000100;
		if(({row_reg, col_reg}==12'b010110011110)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}>=12'b010110011111) && ({row_reg, col_reg}<12'b010110100001)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b010110100001) && ({row_reg, col_reg}<12'b010111000001)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b010111000001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b010111000010)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010111000011)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b010111000100)) color_data = 12'b101100110111;
		if(({row_reg, col_reg}==12'b010111000101)) color_data = 12'b100101011000;
		if(({row_reg, col_reg}==12'b010111000110)) color_data = 12'b011001101010;
		if(({row_reg, col_reg}==12'b010111000111)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==12'b010111001000)) color_data = 12'b001001011000;
		if(({row_reg, col_reg}==12'b010111001001)) color_data = 12'b001101000110;
		if(({row_reg, col_reg}==12'b010111001010)) color_data = 12'b011100100101;
		if(({row_reg, col_reg}==12'b010111001011)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}>=12'b010111001100) && ({row_reg, col_reg}<12'b010111001110)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010111001110)) color_data = 12'b110000100111;
		if(({row_reg, col_reg}==12'b010111001111)) color_data = 12'b101100110111;
		if(({row_reg, col_reg}==12'b010111010000)) color_data = 12'b100000110101;
		if(({row_reg, col_reg}==12'b010111010001)) color_data = 12'b101000110110;
		if(({row_reg, col_reg}==12'b010111010010)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b010111010011)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b010111010100)) color_data = 12'b100000110111;
		if(({row_reg, col_reg}==12'b010111010101)) color_data = 12'b011001011000;
		if(({row_reg, col_reg}==12'b010111010110)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==12'b010111010111)) color_data = 12'b001101101010;
		if(({row_reg, col_reg}==12'b010111011000)) color_data = 12'b011001001000;
		if(({row_reg, col_reg}==12'b010111011001)) color_data = 12'b101000110111;
		if(({row_reg, col_reg}==12'b010111011010)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010111011011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b010111011100)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b010111011101)) color_data = 12'b110100100101;
		if(({row_reg, col_reg}==12'b010111011110)) color_data = 12'b110100010101;
		if(({row_reg, col_reg}==12'b010111011111)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b010111100000) && ({row_reg, col_reg}<12'b011000000001)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011000000001)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b011000000010)) color_data = 12'b110000110111;
		if(({row_reg, col_reg}==12'b011000000011)) color_data = 12'b101001001000;
		if(({row_reg, col_reg}==12'b011000000100)) color_data = 12'b100001111010;
		if(({row_reg, col_reg}==12'b011000000101)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==12'b011000000110)) color_data = 12'b001101101010;
		if(({row_reg, col_reg}==12'b011000000111)) color_data = 12'b001101011000;
		if(({row_reg, col_reg}==12'b011000001000)) color_data = 12'b010001101000;
		if(({row_reg, col_reg}==12'b011000001001)) color_data = 12'b011101101000;
		if(({row_reg, col_reg}==12'b011000001010)) color_data = 12'b101101011000;
		if(({row_reg, col_reg}==12'b011000001011)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b011000001100)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b011000001101)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b011000001110)) color_data = 12'b100101001000;
		if(({row_reg, col_reg}==12'b011000001111)) color_data = 12'b011101001000;
		if(({row_reg, col_reg}==12'b011000010000)) color_data = 12'b011000110101;
		if(({row_reg, col_reg}==12'b011000010001)) color_data = 12'b100001000111;
		if(({row_reg, col_reg}==12'b011000010010)) color_data = 12'b100101000111;
		if(({row_reg, col_reg}==12'b011000010011)) color_data = 12'b100001001000;
		if(({row_reg, col_reg}==12'b011000010100)) color_data = 12'b010001011000;
		if(({row_reg, col_reg}==12'b011000010101)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==12'b011000010110)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==12'b011000010111)) color_data = 12'b001101101001;
		if(({row_reg, col_reg}==12'b011000011000)) color_data = 12'b011101011000;
		if(({row_reg, col_reg}==12'b011000011001)) color_data = 12'b101001000111;
		if(({row_reg, col_reg}==12'b011000011010)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b011000011011)) color_data = 12'b111100010101;
		if(({row_reg, col_reg}==12'b011000011100)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}>=12'b011000011101) && ({row_reg, col_reg}<12'b011000011111)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011000011111)) color_data = 12'b111000010101;

		if(({row_reg, col_reg}>=12'b011000100000) && ({row_reg, col_reg}<12'b011001000000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011001000000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011001000001)) color_data = 12'b110100010110;
		if(({row_reg, col_reg}==12'b011001000010)) color_data = 12'b110000110111;
		if(({row_reg, col_reg}==12'b011001000011)) color_data = 12'b101101011001;
		if(({row_reg, col_reg}==12'b011001000100)) color_data = 12'b100001111011;
		if(({row_reg, col_reg}==12'b011001000101)) color_data = 12'b011001111010;
		if(({row_reg, col_reg}==12'b011001000110)) color_data = 12'b011101111011;
		if(({row_reg, col_reg}==12'b011001000111)) color_data = 12'b100110001100;
		if(({row_reg, col_reg}==12'b011001001000)) color_data = 12'b101010001011;
		if(({row_reg, col_reg}==12'b011001001001)) color_data = 12'b101101101001;
		if(({row_reg, col_reg}==12'b011001001010)) color_data = 12'b110001001000;
		if(({row_reg, col_reg}==12'b011001001011)) color_data = 12'b101100100110;
		if(({row_reg, col_reg}==12'b011001001100)) color_data = 12'b101100110111;
		if(({row_reg, col_reg}==12'b011001001101)) color_data = 12'b100101001000;
		if(({row_reg, col_reg}==12'b011001001110)) color_data = 12'b011001011001;
		if(({row_reg, col_reg}==12'b011001001111)) color_data = 12'b010101101001;
		if(({row_reg, col_reg}==12'b011001010000)) color_data = 12'b010001000111;
		if(({row_reg, col_reg}==12'b011001010001)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==12'b011001010010)) color_data = 12'b100001000111;
		if(({row_reg, col_reg}==12'b011001010011)) color_data = 12'b011101000111;
		if(({row_reg, col_reg}==12'b011001010100)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==12'b011001010101)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==12'b011001010110)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==12'b011001010111)) color_data = 12'b100110001100;
		if(({row_reg, col_reg}==12'b011001011000)) color_data = 12'b110110011100;
		if(({row_reg, col_reg}==12'b011001011001)) color_data = 12'b110101001000;
		if(({row_reg, col_reg}==12'b011001011010)) color_data = 12'b110100010101;
		if(({row_reg, col_reg}==12'b011001011011)) color_data = 12'b111100010101;
		if(({row_reg, col_reg}==12'b011001011100)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}==12'b011001011101)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011001011110)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b011001011111)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b011001100000) && ({row_reg, col_reg}<12'b011010000000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011010000000)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}>=12'b011010000001) && ({row_reg, col_reg}<12'b011010000011)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011010000011)) color_data = 12'b110100110111;
		if(({row_reg, col_reg}==12'b011010000100)) color_data = 12'b110101011001;
		if(({row_reg, col_reg}==12'b011010000101)) color_data = 12'b110101101010;
		if(({row_reg, col_reg}==12'b011010000110)) color_data = 12'b110101011001;
		if(({row_reg, col_reg}==12'b011010000111)) color_data = 12'b110000110111;
		if(({row_reg, col_reg}==12'b011010001000)) color_data = 12'b101100100111;
		if(({row_reg, col_reg}==12'b011010001001)) color_data = 12'b101100100110;
		if(({row_reg, col_reg}==12'b011010001010)) color_data = 12'b101100110111;
		if(({row_reg, col_reg}==12'b011010001011)) color_data = 12'b100101001000;
		if(({row_reg, col_reg}==12'b011010001100)) color_data = 12'b011001011001;
		if(({row_reg, col_reg}==12'b011010001101)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}==12'b011010001110)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==12'b011010001111)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==12'b011010010000)) color_data = 12'b001001101001;
		if(({row_reg, col_reg}==12'b011010010001)) color_data = 12'b010101011000;
		if(({row_reg, col_reg}==12'b011010010010)) color_data = 12'b100100110111;
		if(({row_reg, col_reg}==12'b011010010011)) color_data = 12'b101101001000;
		if(({row_reg, col_reg}==12'b011010010100)) color_data = 12'b101101101001;
		if(({row_reg, col_reg}==12'b011010010101)) color_data = 12'b101001101000;
		if(({row_reg, col_reg}==12'b011010010110)) color_data = 12'b110001101010;
		if(({row_reg, col_reg}==12'b011010010111)) color_data = 12'b110001011001;
		if(({row_reg, col_reg}==12'b011010011000)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}>=12'b011010011001) && ({row_reg, col_reg}<12'b011010011011)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b011010011011)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}==12'b011010011100)) color_data = 12'b111000010101;

		if(({row_reg, col_reg}>=12'b011010011101) && ({row_reg, col_reg}<12'b011011000000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011011000000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011011000001)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}>=12'b011011000010) && ({row_reg, col_reg}<12'b011011000100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011011000100)) color_data = 12'b110100100101;
		if(({row_reg, col_reg}>=12'b011011000101) && ({row_reg, col_reg}<12'b011011000111)) color_data = 12'b110100010101;
		if(({row_reg, col_reg}>=12'b011011000111) && ({row_reg, col_reg}<12'b011011001001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011011001001)) color_data = 12'b110100100111;
		if(({row_reg, col_reg}==12'b011011001010)) color_data = 12'b101001001000;
		if(({row_reg, col_reg}==12'b011011001011)) color_data = 12'b100001101001;
		if(({row_reg, col_reg}==12'b011011001100)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==12'b011011001101)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}==12'b011011001110)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==12'b011011001111)) color_data = 12'b001001011001;
		if(({row_reg, col_reg}==12'b011011010000)) color_data = 12'b001001011000;
		if(({row_reg, col_reg}==12'b011011010001)) color_data = 12'b011001011001;
		if(({row_reg, col_reg}==12'b011011010010)) color_data = 12'b101100111000;
		if(({row_reg, col_reg}==12'b011011010011)) color_data = 12'b110100100111;
		if(({row_reg, col_reg}>=12'b011011010100) && ({row_reg, col_reg}<12'b011011010110)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b011011010110)) color_data = 12'b110000100110;
		if(({row_reg, col_reg}==12'b011011010111)) color_data = 12'b110100010101;
		if(({row_reg, col_reg}>=12'b011011011000) && ({row_reg, col_reg}<12'b011011011011)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011011011011)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}==12'b011011011100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011011011101)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}==12'b011011011110)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b011011011111) && ({row_reg, col_reg}<12'b011100000000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011100000000)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}>=12'b011100000001) && ({row_reg, col_reg}<12'b011100000110)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b011100000110) && ({row_reg, col_reg}<12'b011100001000)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}==12'b011100001000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011100001001)) color_data = 12'b101100100110;
		if(({row_reg, col_reg}==12'b011100001010)) color_data = 12'b011101000111;
		if(({row_reg, col_reg}==12'b011100001011)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==12'b011100001100)) color_data = 12'b001101101001;
		if(({row_reg, col_reg}==12'b011100001101)) color_data = 12'b001001101001;
		if(({row_reg, col_reg}==12'b011100001110)) color_data = 12'b001101101001;
		if(({row_reg, col_reg}==12'b011100001111)) color_data = 12'b011101111010;
		if(({row_reg, col_reg}==12'b011100010000)) color_data = 12'b101110001011;
		if(({row_reg, col_reg}==12'b011100010001)) color_data = 12'b110110001011;
		if(({row_reg, col_reg}==12'b011100010010)) color_data = 12'b110100110111;
		if(({row_reg, col_reg}==12'b011100010011)) color_data = 12'b110100010110;
		if(({row_reg, col_reg}==12'b011100010100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011100010101)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}>=12'b011100010110) && ({row_reg, col_reg}<12'b011100011000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b011100011000) && ({row_reg, col_reg}<12'b011100011010)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b011100011010)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}==12'b011100011011)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b011100011100) && ({row_reg, col_reg}<12'b011100011111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011100011111)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b011100100000) && ({row_reg, col_reg}<12'b011101000000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b011101000000) && ({row_reg, col_reg}<12'b011101000010)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b011101000010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b011101000011) && ({row_reg, col_reg}<12'b011101000110)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011101000110)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}>=12'b011101000111) && ({row_reg, col_reg}<12'b011101001001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011101001001)) color_data = 12'b101100100110;
		if(({row_reg, col_reg}==12'b011101001010)) color_data = 12'b100001001000;
		if(({row_reg, col_reg}==12'b011101001011)) color_data = 12'b100001101010;
		if(({row_reg, col_reg}==12'b011101001100)) color_data = 12'b011101101010;
		if(({row_reg, col_reg}==12'b011101001101)) color_data = 12'b100001111010;
		if(({row_reg, col_reg}==12'b011101001110)) color_data = 12'b101001111011;
		if(({row_reg, col_reg}==12'b011101001111)) color_data = 12'b101101111010;
		if(({row_reg, col_reg}==12'b011101010000)) color_data = 12'b101101000111;
		if(({row_reg, col_reg}==12'b011101010001)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==12'b011101010010)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}>=12'b011101010011) && ({row_reg, col_reg}<12'b011101010111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b011101010111) && ({row_reg, col_reg}<12'b011101011001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011101011001)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}>=12'b011101011010) && ({row_reg, col_reg}<12'b011101011100)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b011101011100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b011101011101) && ({row_reg, col_reg}<12'b011101011111)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b011101011111) && ({row_reg, col_reg}<12'b011110000000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011110000000)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b011110000001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b011110000010) && ({row_reg, col_reg}<12'b011110000101)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011110000101)) color_data = 12'b111100010110;
		if(({row_reg, col_reg}>=12'b011110000110) && ({row_reg, col_reg}<12'b011110001000)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b011110001000)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}==12'b011110001001)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011110001010)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==12'b011110001011)) color_data = 12'b110100110111;
		if(({row_reg, col_reg}==12'b011110001100)) color_data = 12'b110101001000;
		if(({row_reg, col_reg}==12'b011110001101)) color_data = 12'b110001001000;
		if(({row_reg, col_reg}==12'b011110001110)) color_data = 12'b101100100110;
		if(({row_reg, col_reg}>=12'b011110001111) && ({row_reg, col_reg}<12'b011110010001)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==12'b011110010001)) color_data = 12'b110100100101;
		if(({row_reg, col_reg}==12'b011110010010)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b011110010011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011110010100)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011110010101)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011110010110)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}>=12'b011110010111) && ({row_reg, col_reg}<12'b011110011011)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b011110011011) && ({row_reg, col_reg}<12'b011110011101)) color_data = 12'b111000100110;

		if(({row_reg, col_reg}>=12'b011110011101) && ({row_reg, col_reg}<12'b011111000111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011111000111)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b011111001000) && ({row_reg, col_reg}<12'b011111001010)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}>=12'b011111001010) && ({row_reg, col_reg}<12'b011111001100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}>=12'b011111001100) && ({row_reg, col_reg}<12'b011111001110)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}>=12'b011111001110) && ({row_reg, col_reg}<12'b011111010001)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}==12'b011111010001)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b011111010010)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}>=12'b011111010011) && ({row_reg, col_reg}<12'b011111010101)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b011111010101)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011111010110)) color_data = 12'b111100010110;
		if(({row_reg, col_reg}>=12'b011111010111) && ({row_reg, col_reg}<12'b011111011100)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b011111011100)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b011111011101)) color_data = 12'b111000100101;
		if(({row_reg, col_reg}==12'b011111011110)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==12'b011111011111)) color_data = 12'b111000010101;

		if(({row_reg, col_reg}>=12'b011111100000) && ({row_reg, col_reg}<12'b100000001000)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b100000001000)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=12'b100000001001) && ({row_reg, col_reg}<12'b100000001111)) color_data = 12'b111000010110;
		if(({row_reg, col_reg}==12'b100000001111)) color_data = 12'b111000010101;
		if(({row_reg, col_reg}==12'b100000010000)) color_data = 12'b111000100110;





		if(({row_reg, col_reg}>=12'b100000010001) && ({row_reg, col_reg}<=12'b100100100100)) color_data = 12'b111000010110;
	end
endmodule