module gandhi_down_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=12'b000000000000) && ({row_reg, col_reg}<12'b000000010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000000010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b000000010110) && ({row_reg, col_reg}<12'b000000011100)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b000000011100) && ({row_reg, col_reg}<12'b000001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000001010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b000001010100) && ({row_reg, col_reg}<12'b000001011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000001011110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b000001011111) && ({row_reg, col_reg}<12'b000010010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000010010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b000010010010) && ({row_reg, col_reg}<12'b000010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b000010010100) && ({row_reg, col_reg}<12'b000010011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000010011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b000010011101) && ({row_reg, col_reg}<12'b000010011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000010011111)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b000010100000) && ({row_reg, col_reg}<12'b000011001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000011001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b000011010000) && ({row_reg, col_reg}<12'b000011010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000011010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b000011010011) && ({row_reg, col_reg}<12'b000011010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b000011010101) && ({row_reg, col_reg}<12'b000011010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b000011010111) && ({row_reg, col_reg}<12'b000011011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b000011011010) && ({row_reg, col_reg}<12'b000011011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b000011011100) && ({row_reg, col_reg}<12'b000011011111)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b000011011111) && ({row_reg, col_reg}<12'b000100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000100001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b000100010000) && ({row_reg, col_reg}<12'b000100010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000100010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b000100010100) && ({row_reg, col_reg}<12'b000100010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b000100010110) && ({row_reg, col_reg}<12'b000100011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b000100011010) && ({row_reg, col_reg}<12'b000100011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000100011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b000100011110) && ({row_reg, col_reg}<12'b000100100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000100100001)) color_data = 12'b010001000100;

		if(({row_reg, col_reg}>=12'b000100100010) && ({row_reg, col_reg}<12'b000101001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000101001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000101001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000101001111)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==12'b000101010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000101010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b000101010010) && ({row_reg, col_reg}<12'b000101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b000101010100) && ({row_reg, col_reg}<12'b000101011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000101011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b000101011010) && ({row_reg, col_reg}<12'b000101011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000101011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000101011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b000101011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000101100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000101100010)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b000101100011) && ({row_reg, col_reg}<12'b000110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000110001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000110001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000110001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b000110001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b000110010000) && ({row_reg, col_reg}<12'b000110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b000110010011) && ({row_reg, col_reg}<12'b000110011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000110011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b000110011010) && ({row_reg, col_reg}<12'b000110011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000110011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000110011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000110011111)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}>=12'b000110100000) && ({row_reg, col_reg}<12'b000110100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b000110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000110100011)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b000110100100) && ({row_reg, col_reg}<12'b000111001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000111001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000111001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000111001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b000111001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b000111001111) && ({row_reg, col_reg}<12'b000111010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b000111010010) && ({row_reg, col_reg}<12'b000111010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000111010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b000111010110) && ({row_reg, col_reg}<12'b000111011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000111011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000111011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b000111011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000111011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000111011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000111011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b000111011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b000111100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b000111100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b000111100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b000111100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b000111100100)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b000111100101) && ({row_reg, col_reg}<12'b001000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001000001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001000001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001000001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001000001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001000010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001000010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b001000010010) && ({row_reg, col_reg}<12'b001000010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b001000010100) && ({row_reg, col_reg}<12'b001000010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001000010110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=12'b001000010111) && ({row_reg, col_reg}<12'b001000011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001000011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001000011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b001000011111) && ({row_reg, col_reg}<12'b001000100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001000100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001000100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001000100011)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=12'b001000100100) && ({row_reg, col_reg}<12'b001001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001001001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001001001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001001001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001001001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001001001110)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}>=12'b001001001111) && ({row_reg, col_reg}<12'b001001010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001001010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b001001010100) && ({row_reg, col_reg}<12'b001001011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b001001011001) && ({row_reg, col_reg}<12'b001001011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001001011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001001011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001001011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001001011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001001100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b001001100001) && ({row_reg, col_reg}<12'b001001100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001001100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001001100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001001100101)) color_data = 12'b010001000100;

		if(({row_reg, col_reg}>=12'b001001100110) && ({row_reg, col_reg}<12'b001010001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001010001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001010001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001010001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b001010001110) && ({row_reg, col_reg}<12'b001010010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001010010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b001010010001) && ({row_reg, col_reg}<12'b001010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001010011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b001010011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001010100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001010100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001010100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001010100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001010100100)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b001010100101) && ({row_reg, col_reg}<12'b001011001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001011001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001011001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001011001011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001011001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001011001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b001011001110) && ({row_reg, col_reg}<12'b001011010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001011010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b001011010010) && ({row_reg, col_reg}<12'b001011010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001011010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b001011010101) && ({row_reg, col_reg}<12'b001011011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001011011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001011100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001011100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b001011100010) && ({row_reg, col_reg}<12'b001011100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001011100100)) color_data = 12'b010001000100;

		if(({row_reg, col_reg}>=12'b001011100101) && ({row_reg, col_reg}<12'b001100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001100001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b001100001011) && ({row_reg, col_reg}<12'b001100001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b001100010000) && ({row_reg, col_reg}<12'b001100011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001100011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b001100100001) && ({row_reg, col_reg}<12'b001100100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001100100011)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==12'b001100100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001100100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001100100110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b001100100111) && ({row_reg, col_reg}<12'b001101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001101001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001101001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b001101001011) && ({row_reg, col_reg}<12'b001101001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001101001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b001101001110) && ({row_reg, col_reg}<12'b001101010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b001101010000) && ({row_reg, col_reg}<12'b001101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001101011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001101100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001101100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001101100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b001101100011) && ({row_reg, col_reg}<12'b001101100101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001101100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001101100110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b001101100111) && ({row_reg, col_reg}<12'b001110001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001110001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001110001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b001110001011) && ({row_reg, col_reg}<12'b001110001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001110001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001110001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001110001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001110010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b001110010001) && ({row_reg, col_reg}<12'b001110011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001110011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001110100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001110100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001110100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001110100100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001110100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001110100110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b001110100111) && ({row_reg, col_reg}<12'b001111001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001111001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001111001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001111001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001111001100)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b001111001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001111001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001111010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b001111010001) && ({row_reg, col_reg}<12'b001111100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001111100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b001111100001) && ({row_reg, col_reg}<12'b001111100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001111100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001111100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b001111100101) && ({row_reg, col_reg}<12'b001111100111)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b001111100111) && ({row_reg, col_reg}<12'b010000001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010000001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010000001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b010000001011) && ({row_reg, col_reg}<12'b010000001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010000001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010000010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b010000010001) && ({row_reg, col_reg}<12'b010000010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b010000010111) && ({row_reg, col_reg}<12'b010000011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010000011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b010000011010) && ({row_reg, col_reg}<12'b010000100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010000100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010000100001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010000100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010000100011) && ({row_reg, col_reg}<12'b010000100101)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b010000100101) && ({row_reg, col_reg}<12'b010001001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010001001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010001001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010001001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010001001100) && ({row_reg, col_reg}<12'b010001001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010001001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b010001001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b010001010000) && ({row_reg, col_reg}<12'b010001010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010001010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b010001010100) && ({row_reg, col_reg}<12'b010001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010001010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b010001011000) && ({row_reg, col_reg}<12'b010001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b010001011010) && ({row_reg, col_reg}<12'b010001100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010001100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010001100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010001100011) && ({row_reg, col_reg}<12'b010001100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010001100110)) color_data = 12'b011101110101;

		if(({row_reg, col_reg}>=12'b010001100111) && ({row_reg, col_reg}<12'b010010001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010010001001)) color_data = 12'b111111110000;
		if(({row_reg, col_reg}==12'b010010001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010010001011) && ({row_reg, col_reg}<12'b010010001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010010001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010010001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=12'b010010010000) && ({row_reg, col_reg}<12'b010010010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010010010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010010010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b010010010111) && ({row_reg, col_reg}<12'b010010011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b010010011100) && ({row_reg, col_reg}<12'b010010011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010010011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010010011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010010100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010010100010)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==12'b010010100011)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}>=12'b010010100100) && ({row_reg, col_reg}<12'b010010100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010010100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010010101000)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b010010101001) && ({row_reg, col_reg}<12'b010011001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b010011001010) && ({row_reg, col_reg}<12'b010011001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010011001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010011001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010011001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b010011010000) && ({row_reg, col_reg}<12'b010011010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010011010100)) color_data = 12'b100101100110;
		if(({row_reg, col_reg}==12'b010011010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b010011010110) && ({row_reg, col_reg}<12'b010011011000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010011011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010011011001) && ({row_reg, col_reg}<12'b010011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010011011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b010011011111) && ({row_reg, col_reg}<12'b010011100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b010011100001) && ({row_reg, col_reg}<12'b010011100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b010011100011) && ({row_reg, col_reg}<12'b010011100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010011100101)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==12'b010011100110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010011101000)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b010011101001) && ({row_reg, col_reg}<12'b010100001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010100001000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010100001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010100001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010100001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b010100001100) && ({row_reg, col_reg}<12'b010100001110)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==12'b010100001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010100010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b010100010001) && ({row_reg, col_reg}<12'b010100010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010100010100)) color_data = 12'b111011101100;
		if(({row_reg, col_reg}==12'b010100010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010100010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010100010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b010100011000) && ({row_reg, col_reg}<12'b010100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010100011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010100011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b010100011110) && ({row_reg, col_reg}<12'b010100100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010100100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b010100100001) && ({row_reg, col_reg}<12'b010100100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010100100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010100100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b010100100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010100100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010100100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010100101000)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b010100101001) && ({row_reg, col_reg}<12'b010101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010101001000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010101001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010101001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010101001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010101001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010101001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010101001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010101001111) && ({row_reg, col_reg}<12'b010101010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010101010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010101010100) && ({row_reg, col_reg}<12'b010101010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010101010111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==12'b010101011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010101011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b010101011010) && ({row_reg, col_reg}<12'b010101011100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}>=12'b010101011100) && ({row_reg, col_reg}<12'b010101011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010101011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010101011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010101100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b010101100001) && ({row_reg, col_reg}<12'b010101100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010101100011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010101100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b010101100101) && ({row_reg, col_reg}<12'b010101100111)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b010101100111) && ({row_reg, col_reg}<12'b010110001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b010110001010) && ({row_reg, col_reg}<12'b010110001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010110001100) && ({row_reg, col_reg}<12'b010110001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010110001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010110001111) && ({row_reg, col_reg}<12'b010110010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b010110010001) && ({row_reg, col_reg}<12'b010110010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010110010011) && ({row_reg, col_reg}<12'b010110010101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b010110010101) && ({row_reg, col_reg}<12'b010110011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010110011001) && ({row_reg, col_reg}<12'b010110011011)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}>=12'b010110011011) && ({row_reg, col_reg}<12'b010110011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010110011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010110011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010110100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010110100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b010110100010) && ({row_reg, col_reg}<12'b010110100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010110100101)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b010110100110) && ({row_reg, col_reg}<12'b010111001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010111001001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010111001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010111001101)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==12'b010111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010111001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111010000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010111010001)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b010111010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010111010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b010111010100) && ({row_reg, col_reg}<12'b010111011000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010111011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b010111011010) && ({row_reg, col_reg}<12'b010111011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111011100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010111011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111011110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b010111011111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010111100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010111100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010111100011)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==12'b010111100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010111100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010111100111)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b010111101000) && ({row_reg, col_reg}<12'b011000001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011000001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011000001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011000001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011000001100)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==12'b011000001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b011000001110) && ({row_reg, col_reg}<12'b011000010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011000010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011000010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011000010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011000010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011000010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011000011000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011000011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011000011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011000011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011000011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011000011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011000100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011000100001)) color_data = 12'b011001010110;
		if(({row_reg, col_reg}==12'b011000100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011000100011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==12'b011000100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000100101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011000100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011000100111)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b011000101000) && ({row_reg, col_reg}<12'b011001001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011001001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b011001001100) && ({row_reg, col_reg}<12'b011001001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011001001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b011001001111) && ({row_reg, col_reg}<12'b011001010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011001010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011001010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011001010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011001011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011001011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011001011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011001011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=12'b011001011100) && ({row_reg, col_reg}<12'b011001011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011001011110) && ({row_reg, col_reg}<12'b011001100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011001100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011001100001) && ({row_reg, col_reg}<12'b011001100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011001100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011001100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011001100101)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=12'b011001100110) && ({row_reg, col_reg}<12'b011010001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011010001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011010001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011010001100) && ({row_reg, col_reg}<12'b011010001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011010001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b011010001111) && ({row_reg, col_reg}<12'b011010010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011010010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b011010010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011010010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=12'b011010011000) && ({row_reg, col_reg}<12'b011010011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011010011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b011010011100) && ({row_reg, col_reg}<12'b011010100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011010100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011010100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011010100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011010100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011010100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011010100101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011010100110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b011010100111) && ({row_reg, col_reg}<12'b011011001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011011001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011011001100) && ({row_reg, col_reg}<12'b011011001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011011001110)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b011011001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b011011010000) && ({row_reg, col_reg}<12'b011011010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011011010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011011010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011011010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011011010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011011011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b011011011001) && ({row_reg, col_reg}<12'b011011011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011011011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011011011111) && ({row_reg, col_reg}<12'b011011100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b011011100001) && ({row_reg, col_reg}<12'b011011100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011011100100)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=12'b011011100101) && ({row_reg, col_reg}<12'b011100001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011100001101) && ({row_reg, col_reg}<12'b011100001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b011100001111) && ({row_reg, col_reg}<12'b011100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011100010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011100010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011100010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011100010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011100010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011100010111) && ({row_reg, col_reg}<12'b011100011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011100011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011100011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b011100011011) && ({row_reg, col_reg}<12'b011100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011100011110) && ({row_reg, col_reg}<12'b011100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011100100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b011100100001) && ({row_reg, col_reg}<12'b011100100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011100100011)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=12'b011100100100) && ({row_reg, col_reg}<12'b011101001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011101001100)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011101001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011101001110) && ({row_reg, col_reg}<12'b011101010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011101010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011101010001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011101010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b011101010011) && ({row_reg, col_reg}<12'b011101010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011101010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011101010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011101010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011101011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011101011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011101011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011101011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011101011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011101011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011101011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b011101100000) && ({row_reg, col_reg}<12'b011101100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b011101100010) && ({row_reg, col_reg}<12'b011101100100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011101100100)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b011101100101) && ({row_reg, col_reg}<12'b011110001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011110001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011110001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b011110001110) && ({row_reg, col_reg}<12'b011110010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011110010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011110010011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b011110010100) && ({row_reg, col_reg}<12'b011110010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011110010111) && ({row_reg, col_reg}<12'b011110011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011110011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011110011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011110011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b011110011101) && ({row_reg, col_reg}<12'b011110100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011110100000) && ({row_reg, col_reg}<12'b011110100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b011110100011) && ({row_reg, col_reg}<12'b011110100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b011110100110) && ({row_reg, col_reg}<12'b011110101000)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b011110101000) && ({row_reg, col_reg}<12'b011111001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011111001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b011111001100) && ({row_reg, col_reg}<12'b011111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011111001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011111001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011111010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011111010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011111010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011111010011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011111010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b011111010101) && ({row_reg, col_reg}<12'b011111011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b011111011000) && ({row_reg, col_reg}<12'b011111011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011111011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b011111011100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b011111011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011111011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011111011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011111100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011111100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011111100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011111100011)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}>=12'b011111100100) && ({row_reg, col_reg}<12'b011111100110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b011111100110) && ({row_reg, col_reg}<12'b011111101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b011111101001)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b011111101010) && ({row_reg, col_reg}<12'b100000001001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100000001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100000001010) && ({row_reg, col_reg}<12'b100000001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100000001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100000001101) && ({row_reg, col_reg}<12'b100000010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100000010000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b100000010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100000010010) && ({row_reg, col_reg}<12'b100000010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100000010100) && ({row_reg, col_reg}<12'b100000010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100000010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100000010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100000011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100000011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100000011010) && ({row_reg, col_reg}<12'b100000011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100000011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100000011101)) color_data = 12'b010001001000;
		if(({row_reg, col_reg}==12'b100000011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100000011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100000100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100000100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100000100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100000100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100000100100) && ({row_reg, col_reg}<12'b100000101000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100000101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b100000101001) && ({row_reg, col_reg}<12'b100000101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100000101011)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b100000101100) && ({row_reg, col_reg}<12'b100001000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100001000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100001001000) && ({row_reg, col_reg}<12'b100001001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100001001010) && ({row_reg, col_reg}<12'b100001001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100001001111) && ({row_reg, col_reg}<12'b100001010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100001010010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001010011)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b100001010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100001010110) && ({row_reg, col_reg}<12'b100001011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100001011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100001011111) && ({row_reg, col_reg}<12'b100001100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100001100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100001100100) && ({row_reg, col_reg}<12'b100001100110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100001100110) && ({row_reg, col_reg}<12'b100001101011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100001101011) && ({row_reg, col_reg}<12'b100001101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100001101101)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b100001101110) && ({row_reg, col_reg}<12'b100010000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100010000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b100010000101) && ({row_reg, col_reg}<12'b100010001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100010001000) && ({row_reg, col_reg}<12'b100010001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100010001100) && ({row_reg, col_reg}<12'b100010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100010001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b100010001111) && ({row_reg, col_reg}<12'b100010010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100010010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100010010010) && ({row_reg, col_reg}<12'b100010010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100010010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100010010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100010010110) && ({row_reg, col_reg}<12'b100010011000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100010011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100010011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=12'b100010011010) && ({row_reg, col_reg}<12'b100010011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100010011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100010011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100010011110) && ({row_reg, col_reg}<12'b100010100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100010100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100010100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100010100010) && ({row_reg, col_reg}<12'b100010100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100010100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100010100101) && ({row_reg, col_reg}<12'b100010101000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100010101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100010101001) && ({row_reg, col_reg}<12'b100010101101)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b100010101101) && ({row_reg, col_reg}<12'b100011000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100011000110) && ({row_reg, col_reg}<12'b100011001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100011001010) && ({row_reg, col_reg}<12'b100011001101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100011001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100011001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100011001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100011010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100011010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100011010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100011010011) && ({row_reg, col_reg}<12'b100011010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b100011010101) && ({row_reg, col_reg}<12'b100011010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100011010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100011011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100011011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100011011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100011011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100011011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100011011101) && ({row_reg, col_reg}<12'b100011100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100011100000) && ({row_reg, col_reg}<12'b100011100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100011100010) && ({row_reg, col_reg}<12'b100011100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100011100100) && ({row_reg, col_reg}<12'b100011100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100011100111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100011101000) && ({row_reg, col_reg}<12'b100011101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100011101011) && ({row_reg, col_reg}<12'b100011101110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100011101110)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=12'b100011101111) && ({row_reg, col_reg}<12'b100100000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100100000100) && ({row_reg, col_reg}<12'b100100001000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100100001000) && ({row_reg, col_reg}<12'b100100001010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100100001010) && ({row_reg, col_reg}<12'b100100001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100100001100) && ({row_reg, col_reg}<12'b100100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100100001110) && ({row_reg, col_reg}<12'b100100010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100100010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100100010001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100100010010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100100010011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==12'b100100010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b100100010101) && ({row_reg, col_reg}<12'b100100010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100100010111)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==12'b100100011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100100011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100100011011) && ({row_reg, col_reg}<12'b100100100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100100100000) && ({row_reg, col_reg}<12'b100100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100100100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100100100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100100100100) && ({row_reg, col_reg}<12'b100100101001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100100101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100100101010) && ({row_reg, col_reg}<12'b100100101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100100101101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100100101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100100101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100100110000)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}==12'b100100110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b100101000000) && ({row_reg, col_reg}<12'b100101000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100101000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100101000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b100101000100) && ({row_reg, col_reg}<12'b100101000110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100101000110) && ({row_reg, col_reg}<12'b100101001000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100101001001) && ({row_reg, col_reg}<12'b100101001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100101001110) && ({row_reg, col_reg}<12'b100101010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100101010000) && ({row_reg, col_reg}<12'b100101010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100101010010) && ({row_reg, col_reg}<12'b100101010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100101010101) && ({row_reg, col_reg}<12'b100101011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100101011010) && ({row_reg, col_reg}<12'b100101011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100101011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100101011101) && ({row_reg, col_reg}<12'b100101011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100101100000)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100101100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100101100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100101100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100101100100) && ({row_reg, col_reg}<12'b100101101011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100101101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100101101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100101101101) && ({row_reg, col_reg}<12'b100101101111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100101101111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=12'b100101110000) && ({row_reg, col_reg}<12'b100110000010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100110000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b100110000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100110000100) && ({row_reg, col_reg}<12'b100110000110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100110000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100110000111) && ({row_reg, col_reg}<12'b100110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100110001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100110001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100110010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100110010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100110010011) && ({row_reg, col_reg}<12'b100110011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100110011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100110011100) && ({row_reg, col_reg}<12'b100110011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100110011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100110011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100110100000) && ({row_reg, col_reg}<12'b100110100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100110100010) && ({row_reg, col_reg}<12'b100110100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100110100100) && ({row_reg, col_reg}<12'b100110101110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100110101110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b100110101111) && ({row_reg, col_reg}<12'b100111000100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100111000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b100111000101) && ({row_reg, col_reg}<12'b100111001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100111001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100111001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100111010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100111010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100111010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b100111010011) && ({row_reg, col_reg}<12'b100111010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100111010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b100111010110) && ({row_reg, col_reg}<12'b100111011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100111011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100111011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b100111011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100111011100)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==12'b100111011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100111011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b100111011111) && ({row_reg, col_reg}<12'b100111100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b100111100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100111100010)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b100111100011) && ({row_reg, col_reg}<12'b101000001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101000001110) && ({row_reg, col_reg}<12'b101000010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101000010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101000010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b101000010010) && ({row_reg, col_reg}<12'b101000010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101000010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101000010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101000010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101000010111) && ({row_reg, col_reg}<12'b101000011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101000011001)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b101000011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101000011011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101000011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b101000011101) && ({row_reg, col_reg}<12'b101000100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101000100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101000100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101000100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101000100100)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b101000100101) && ({row_reg, col_reg}<12'b101001001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101001001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101001001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b101001010000) && ({row_reg, col_reg}<12'b101001010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101001010010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==12'b101001010011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101001010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b101001010101) && ({row_reg, col_reg}<12'b101001010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b101001010111) && ({row_reg, col_reg}<12'b101001011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101001011001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b101001011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101001011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101001011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101001011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b101001011110) && ({row_reg, col_reg}<12'b101001100001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101001100001) && ({row_reg, col_reg}<12'b101001100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101001100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101001100100)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b101001100101) && ({row_reg, col_reg}<12'b101010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101010001110) && ({row_reg, col_reg}<12'b101010010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101010010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101010010001) && ({row_reg, col_reg}<12'b101010010101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101010010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101010010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101010010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101010011000)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b101010011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101010011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b101010011011) && ({row_reg, col_reg}<12'b101010011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101010011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101010100000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101010100001) && ({row_reg, col_reg}<12'b101010100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101010100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101010100100)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b101010100101) && ({row_reg, col_reg}<12'b101011001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101011001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b101011001111) && ({row_reg, col_reg}<12'b101011010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b101011010011) && ({row_reg, col_reg}<12'b101011010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101011010101) && ({row_reg, col_reg}<12'b101011010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b101011010111) && ({row_reg, col_reg}<12'b101011011001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101011011001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b101011011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b101011011011) && ({row_reg, col_reg}<12'b101011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101011011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101011011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b101011100000) && ({row_reg, col_reg}<12'b101011100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101011100010)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}>=12'b101011100011) && ({row_reg, col_reg}<12'b101100001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101100001110) && ({row_reg, col_reg}<12'b101100010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=12'b101100010000) && ({row_reg, col_reg}<12'b101100010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101100010010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101100010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b101100010100) && ({row_reg, col_reg}<12'b101100010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101100010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101100011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b101100011001) && ({row_reg, col_reg}<12'b101100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101100011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101100011100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101100011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101100011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101100011111) && ({row_reg, col_reg}<12'b101100100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101100100010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101100100011)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b101100100100) && ({row_reg, col_reg}<12'b101101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101101001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b101101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b101101010001) && ({row_reg, col_reg}<12'b101101010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101101010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101101010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=12'b101101010110) && ({row_reg, col_reg}<12'b101101011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b101101011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==12'b101101011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b101101011010) && ({row_reg, col_reg}<12'b101101011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101101011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101101011111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101101100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101101100001)) color_data = 12'b010101010101;

		if(({row_reg, col_reg}>=12'b101101100010) && ({row_reg, col_reg}<12'b101110010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101110010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101110010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101110010110) && ({row_reg, col_reg}<12'b101110011000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b101110011000) && ({row_reg, col_reg}<12'b101110011010)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=12'b101110011010) && ({row_reg, col_reg}<12'b101111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b101111010000) && ({row_reg, col_reg}<12'b101111010100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b101111010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==12'b101111010101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=12'b101111010110) && ({row_reg, col_reg}<12'b101111011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b101111011000)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=12'b101111011001) && ({row_reg, col_reg}<12'b110000010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b110000010110)) color_data = 12'b111111111111;


		if(({row_reg, col_reg}>=12'b110000010111) && ({row_reg, col_reg}<=12'b110001110001)) color_data = 12'b000000000000;
	end
endmodule