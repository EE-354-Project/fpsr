module chillguy_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin


		if(({row_reg, col_reg}>=12'b000000000000) && ({row_reg, col_reg}<12'b000010010110)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b000010010110)) color_data = 12'b101000000000;




		if(({row_reg, col_reg}>=12'b000010010111) && ({row_reg, col_reg}<12'b000110011100)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b000110011100) && ({row_reg, col_reg}<12'b000110011110)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b000110011110) && ({row_reg, col_reg}<12'b000111011000)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b000111011000) && ({row_reg, col_reg}<12'b000111011010)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b000111011010) && ({row_reg, col_reg}<12'b000111011110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=12'b000111011110) && ({row_reg, col_reg}<12'b000111100000)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b000111100000) && ({row_reg, col_reg}<12'b001000010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b001000010001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b001000010010) && ({row_reg, col_reg}<12'b001000010111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b001000010111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b001000011000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b001000011001)) color_data = 12'b101000100001;
		if(({row_reg, col_reg}==12'b001000011010)) color_data = 12'b110001010011;
		if(({row_reg, col_reg}==12'b001000011011)) color_data = 12'b011100010000;
		if(({row_reg, col_reg}==12'b001000011100)) color_data = 12'b011100100000;
		if(({row_reg, col_reg}==12'b001000011101)) color_data = 12'b101101010100;
		if(({row_reg, col_reg}==12'b001000011110)) color_data = 12'b101100110010;
		if(({row_reg, col_reg}==12'b001000011111)) color_data = 12'b100100000000;

		if(({row_reg, col_reg}>=12'b001000100000) && ({row_reg, col_reg}<12'b001001010000)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b001001010000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b001001010001) && ({row_reg, col_reg}<12'b001001010111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b001001010111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b001001011000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b001001011001)) color_data = 12'b101101010011;
		if(({row_reg, col_reg}==12'b001001011010)) color_data = 12'b110001110101;
		if(({row_reg, col_reg}==12'b001001011011)) color_data = 12'b011000100000;
		if(({row_reg, col_reg}==12'b001001011100)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==12'b001001011101)) color_data = 12'b101101110101;
		if(({row_reg, col_reg}==12'b001001011110)) color_data = 12'b101101000011;
		if(({row_reg, col_reg}==12'b001001011111)) color_data = 12'b100100000000;

		if(({row_reg, col_reg}>=12'b001001100000) && ({row_reg, col_reg}<12'b001010001011)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b001010001011)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b001010001100) && ({row_reg, col_reg}<12'b001010010111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b001010010111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b001010011000)) color_data = 12'b100100010000;
		if(({row_reg, col_reg}==12'b001010011001)) color_data = 12'b101001000010;
		if(({row_reg, col_reg}==12'b001010011010)) color_data = 12'b101101110101;
		if(({row_reg, col_reg}==12'b001010011011)) color_data = 12'b011000110000;
		if(({row_reg, col_reg}==12'b001010011100)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==12'b001010011101)) color_data = 12'b101001100011;
		if(({row_reg, col_reg}==12'b001010011110)) color_data = 12'b100100100001;
		if(({row_reg, col_reg}==12'b001010011111)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b001010100000) && ({row_reg, col_reg}<12'b001011001001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b001011001001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b001011001010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b001011001011)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b001011001100) && ({row_reg, col_reg}<12'b001011010010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b001011010010) && ({row_reg, col_reg}<12'b001011010101)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b001011010101)) color_data = 12'b101000010000;
		if(({row_reg, col_reg}>=12'b001011010110) && ({row_reg, col_reg}<12'b001011011000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b001011011000)) color_data = 12'b011100010000;
		if(({row_reg, col_reg}==12'b001011011001)) color_data = 12'b100001000010;
		if(({row_reg, col_reg}==12'b001011011010)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==12'b001011011011)) color_data = 12'b011100110001;
		if(({row_reg, col_reg}==12'b001011011100)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==12'b001011011101)) color_data = 12'b100101010010;
		if(({row_reg, col_reg}==12'b001011011110)) color_data = 12'b100100000000;

		if(({row_reg, col_reg}>=12'b001011011111) && ({row_reg, col_reg}<12'b001100001101)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b001100001101)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b001100001110)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b001100001111) && ({row_reg, col_reg}<12'b001100010001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b001100010001)) color_data = 12'b100100010000;
		if(({row_reg, col_reg}==12'b001100010010)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=12'b001100010011) && ({row_reg, col_reg}<12'b001100010101)) color_data = 12'b011100010000;
		if(({row_reg, col_reg}==12'b001100010101)) color_data = 12'b100000100001;
		if(({row_reg, col_reg}==12'b001100010110)) color_data = 12'b100100110010;
		if(({row_reg, col_reg}==12'b001100010111)) color_data = 12'b100101000010;
		if(({row_reg, col_reg}>=12'b001100011000) && ({row_reg, col_reg}<12'b001100011010)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}==12'b001100011010)) color_data = 12'b101001110101;
		if(({row_reg, col_reg}>=12'b001100011011) && ({row_reg, col_reg}<12'b001100011101)) color_data = 12'b101001110100;
		if(({row_reg, col_reg}==12'b001100011101)) color_data = 12'b100000110000;
		if(({row_reg, col_reg}==12'b001100011110)) color_data = 12'b101000010000;

		if(({row_reg, col_reg}>=12'b001100011111) && ({row_reg, col_reg}<12'b001101001001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b001101001001) && ({row_reg, col_reg}<12'b001101001100)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b001101001100)) color_data = 12'b101000010001;
		if(({row_reg, col_reg}>=12'b001101001101) && ({row_reg, col_reg}<12'b001101001111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b001101001111)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==12'b001101010000)) color_data = 12'b100000010000;
		if(({row_reg, col_reg}==12'b001101010001)) color_data = 12'b100000100000;
		if(({row_reg, col_reg}==12'b001101010010)) color_data = 12'b100100110001;
		if(({row_reg, col_reg}==12'b001101010011)) color_data = 12'b101001010011;
		if(({row_reg, col_reg}==12'b001101010100)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==12'b001101010101)) color_data = 12'b011000110000;
		if(({row_reg, col_reg}==12'b001101010110)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==12'b001101010111)) color_data = 12'b101110000101;
		if(({row_reg, col_reg}==12'b001101011000)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==12'b001101011001)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==12'b001101011010)) color_data = 12'b011000110001;
		if(({row_reg, col_reg}==12'b001101011011)) color_data = 12'b101001110100;
		if(({row_reg, col_reg}==12'b001101011100)) color_data = 12'b101110000101;
		if(({row_reg, col_reg}==12'b001101011101)) color_data = 12'b100101000010;
		if(({row_reg, col_reg}==12'b001101011110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b001101011111)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b001101100000) && ({row_reg, col_reg}<12'b001110000111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b001110000111) && ({row_reg, col_reg}<12'b001110001001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b001110001001)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b001110001010)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==12'b001110001011)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==12'b001110001100)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==12'b001110001101)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==12'b001110001110)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}==12'b001110001111)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==12'b001110010000)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}==12'b001110010001)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}>=12'b001110010010) && ({row_reg, col_reg}<12'b001110010100)) color_data = 12'b101110000101;
		if(({row_reg, col_reg}==12'b001110010100)) color_data = 12'b101001110100;
		if(({row_reg, col_reg}==12'b001110010101)) color_data = 12'b011000110001;
		if(({row_reg, col_reg}==12'b001110010110)) color_data = 12'b010000010000;
		if(({row_reg, col_reg}==12'b001110010111)) color_data = 12'b100101110100;
		if(({row_reg, col_reg}==12'b001110011000)) color_data = 12'b100001100011;
		if(({row_reg, col_reg}==12'b001110011001)) color_data = 12'b010100110000;
		if(({row_reg, col_reg}==12'b001110011010)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==12'b001110011011)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==12'b001110011100)) color_data = 12'b100101110100;
		if(({row_reg, col_reg}==12'b001110011101)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==12'b001110011110)) color_data = 12'b100100010000;
		if(({row_reg, col_reg}==12'b001110011111)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b001110100000) && ({row_reg, col_reg}<12'b001111000111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b001111000111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b001111001000)) color_data = 12'b100100000001;
		if(({row_reg, col_reg}==12'b001111001001)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==12'b001111001010)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==12'b001111001011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==12'b001111001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=12'b001111001101) && ({row_reg, col_reg}<12'b001111001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b001111001111)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==12'b001111010000)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}>=12'b001111010001) && ({row_reg, col_reg}<12'b001111010101)) color_data = 12'b101001110100;
		if(({row_reg, col_reg}==12'b001111010101)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==12'b001111010110)) color_data = 12'b010100100000;
		if(({row_reg, col_reg}==12'b001111010111)) color_data = 12'b100101110100;
		if(({row_reg, col_reg}==12'b001111011000)) color_data = 12'b101010010110;
		if(({row_reg, col_reg}==12'b001111011001)) color_data = 12'b010101000001;
		if(({row_reg, col_reg}==12'b001111011010)) color_data = 12'b011101000001;
		if(({row_reg, col_reg}==12'b001111011011)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b001111011100)) color_data = 12'b100110000100;
		if(({row_reg, col_reg}==12'b001111011101)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==12'b001111011110)) color_data = 12'b100100110001;
		if(({row_reg, col_reg}==12'b001111011111)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b001111100000) && ({row_reg, col_reg}<12'b010000000111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b010000000111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b010000001000)) color_data = 12'b100000010000;
		if(({row_reg, col_reg}==12'b010000001001)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}>=12'b010000001010) && ({row_reg, col_reg}<12'b010000001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=12'b010000001100) && ({row_reg, col_reg}<12'b010000001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010000001111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==12'b010000010000)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==12'b010000010001)) color_data = 12'b101001110100;
		if(({row_reg, col_reg}==12'b010000010010)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}>=12'b010000010011) && ({row_reg, col_reg}<12'b010000010101)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}>=12'b010000010101) && ({row_reg, col_reg}<12'b010000011000)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}>=12'b010000011000) && ({row_reg, col_reg}<12'b010000011010)) color_data = 12'b100110000100;
		if(({row_reg, col_reg}>=12'b010000011010) && ({row_reg, col_reg}<12'b010000011100)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b010000011100)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010000011101)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==12'b010000011110)) color_data = 12'b101001000010;
		if(({row_reg, col_reg}==12'b010000011111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b010000100000)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b010000100001) && ({row_reg, col_reg}<12'b010001000111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b010001000111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b010001001000)) color_data = 12'b011100010000;
		if(({row_reg, col_reg}==12'b010001001001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==12'b010001001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=12'b010001001011) && ({row_reg, col_reg}<12'b010001001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010001001111)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==12'b010001010000)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==12'b010001010001)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}>=12'b010001010010) && ({row_reg, col_reg}<12'b010001010101)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010001010101)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}>=12'b010001010110) && ({row_reg, col_reg}<12'b010001011000)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010001011000)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b010001011001)) color_data = 12'b100110000011;
		if(({row_reg, col_reg}==12'b010001011010)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010001011011)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}==12'b010001011100)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010001011101)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==12'b010001011110)) color_data = 12'b101001000010;
		if(({row_reg, col_reg}==12'b010001011111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b010001100000)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b010001100001) && ({row_reg, col_reg}<12'b010010000111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b010010000111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b010010001000)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==12'b010010001001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=12'b010010001010) && ({row_reg, col_reg}<12'b010010001100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010010001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=12'b010010001101) && ({row_reg, col_reg}<12'b010010001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010010001111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==12'b010010010000)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}>=12'b010010010001) && ({row_reg, col_reg}<12'b010010010101)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}>=12'b010010010101) && ({row_reg, col_reg}<12'b010010010111)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}>=12'b010010010111) && ({row_reg, col_reg}<12'b010010011010)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010010011010)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}>=12'b010010011011) && ({row_reg, col_reg}<12'b010010011101)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010010011101)) color_data = 12'b110010000100;
		if(({row_reg, col_reg}==12'b010010011110)) color_data = 12'b101001000010;
		if(({row_reg, col_reg}==12'b010010011111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b010010100000)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b010010100001) && ({row_reg, col_reg}<12'b010011000111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b010011000111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b010011001000)) color_data = 12'b011100010000;
		if(({row_reg, col_reg}==12'b010011001001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==12'b010011001010)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=12'b010011001011) && ({row_reg, col_reg}<12'b010011001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010011001111)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==12'b010011010000)) color_data = 12'b100110000101;
		if(({row_reg, col_reg}>=12'b010011010001) && ({row_reg, col_reg}<12'b010011010011)) color_data = 12'b100110000011;
		if(({row_reg, col_reg}>=12'b010011010011) && ({row_reg, col_reg}<12'b010011010101)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010011010101)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}>=12'b010011010110) && ({row_reg, col_reg}<12'b010011011010)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}>=12'b010011011010) && ({row_reg, col_reg}<12'b010011011100)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b010011011100)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}==12'b010011011101)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==12'b010011011110)) color_data = 12'b101001000010;
		if(({row_reg, col_reg}==12'b010011011111)) color_data = 12'b100100010000;
		if(({row_reg, col_reg}==12'b010011100000)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b010011100001) && ({row_reg, col_reg}<12'b010100000111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b010100000111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b010100001000)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b010100001001)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}>=12'b010100001010) && ({row_reg, col_reg}<12'b010100001100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=12'b010100001100) && ({row_reg, col_reg}<12'b010100001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010100001111)) color_data = 12'b010101010010;
		if(({row_reg, col_reg}==12'b010100010000)) color_data = 12'b100110010101;
		if(({row_reg, col_reg}>=12'b010100010001) && ({row_reg, col_reg}<12'b010100010011)) color_data = 12'b100110000011;
		if(({row_reg, col_reg}==12'b010100010011)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}>=12'b010100010100) && ({row_reg, col_reg}<12'b010100010110)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b010100010110)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010100010111)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}==12'b010100011000)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010100011001)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}>=12'b010100011010) && ({row_reg, col_reg}<12'b010100011100)) color_data = 12'b101001110100;
		if(({row_reg, col_reg}==12'b010100011100)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}==12'b010100011101)) color_data = 12'b110001110101;
		if(({row_reg, col_reg}==12'b010100011110)) color_data = 12'b101101000010;
		if(({row_reg, col_reg}==12'b010100011111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=12'b010100100000) && ({row_reg, col_reg}<12'b010100100010)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b010100100010) && ({row_reg, col_reg}<12'b010101000111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b010101000111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b010101001000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b010101001001)) color_data = 12'b011000000000;
		if(({row_reg, col_reg}==12'b010101001010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==12'b010101001011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=12'b010101001100) && ({row_reg, col_reg}<12'b010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010101001111)) color_data = 12'b011001100011;
		if(({row_reg, col_reg}==12'b010101010000)) color_data = 12'b100110010100;
		if(({row_reg, col_reg}==12'b010101010001)) color_data = 12'b100110000011;
		if(({row_reg, col_reg}>=12'b010101010010) && ({row_reg, col_reg}<12'b010101010100)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010101010100)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}>=12'b010101010101) && ({row_reg, col_reg}<12'b010101011001)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}>=12'b010101011001) && ({row_reg, col_reg}<12'b010101011101)) color_data = 12'b101001110100;
		if(({row_reg, col_reg}==12'b010101011101)) color_data = 12'b110001110100;
		if(({row_reg, col_reg}==12'b010101011110)) color_data = 12'b101000110010;
		if(({row_reg, col_reg}==12'b010101011111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b010101100000)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b010101100001) && ({row_reg, col_reg}<12'b010110001000)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b010110001000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b010110001001)) color_data = 12'b101000000001;
		if(({row_reg, col_reg}==12'b010110001010)) color_data = 12'b010100000000;
		if(({row_reg, col_reg}==12'b010110001011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=12'b010110001100) && ({row_reg, col_reg}<12'b010110001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==12'b010110001110)) color_data = 12'b001000100000;
		if(({row_reg, col_reg}==12'b010110001111)) color_data = 12'b100010000101;
		if(({row_reg, col_reg}==12'b010110010000)) color_data = 12'b100110000100;
		if(({row_reg, col_reg}==12'b010110010001)) color_data = 12'b100110000011;
		if(({row_reg, col_reg}>=12'b010110010010) && ({row_reg, col_reg}<12'b010110010100)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==12'b010110010100)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}>=12'b010110010101) && ({row_reg, col_reg}<12'b010110011001)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b010110011001)) color_data = 12'b100001100010;
		if(({row_reg, col_reg}==12'b010110011010)) color_data = 12'b011101010001;
		if(({row_reg, col_reg}==12'b010110011011)) color_data = 12'b100101110011;
		if(({row_reg, col_reg}==12'b010110011100)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b010110011101)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==12'b010110011110)) color_data = 12'b101000110010;
		if(({row_reg, col_reg}>=12'b010110011111) && ({row_reg, col_reg}<12'b010110100001)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b010110100001) && ({row_reg, col_reg}<12'b010111001001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b010111001001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b010111001010)) color_data = 12'b100100010001;
		if(({row_reg, col_reg}==12'b010111001011)) color_data = 12'b011100010001;
		if(({row_reg, col_reg}==12'b010111001100)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==12'b010111001101)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==12'b010111001110)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}>=12'b010111001111) && ({row_reg, col_reg}<12'b010111010001)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==12'b010111010001)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}>=12'b010111010010) && ({row_reg, col_reg}<12'b010111010100)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}>=12'b010111010100) && ({row_reg, col_reg}<12'b010111010110)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b010111010110)) color_data = 12'b100101110011;
		if(({row_reg, col_reg}==12'b010111010111)) color_data = 12'b100001100010;
		if(({row_reg, col_reg}==12'b010111011000)) color_data = 12'b011101000001;
		if(({row_reg, col_reg}==12'b010111011001)) color_data = 12'b100001010010;
		if(({row_reg, col_reg}==12'b010111011010)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==12'b010111011011)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b010111011100)) color_data = 12'b100101110100;
		if(({row_reg, col_reg}==12'b010111011101)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==12'b010111011110)) color_data = 12'b101000110010;
		if(({row_reg, col_reg}==12'b010111011111)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b010111100000) && ({row_reg, col_reg}<12'b011000001010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b011000001010) && ({row_reg, col_reg}<12'b011000001100)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b011000001100)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==12'b011000001101)) color_data = 12'b100000010000;
		if(({row_reg, col_reg}==12'b011000001110)) color_data = 12'b100000100001;
		if(({row_reg, col_reg}==12'b011000001111)) color_data = 12'b100000110001;
		if(({row_reg, col_reg}==12'b011000010000)) color_data = 12'b100101000001;
		if(({row_reg, col_reg}==12'b011000010001)) color_data = 12'b100101100010;
		if(({row_reg, col_reg}==12'b011000010010)) color_data = 12'b100101110011;
		if(({row_reg, col_reg}==12'b011000010011)) color_data = 12'b100110000011;
		if(({row_reg, col_reg}==12'b011000010100)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b011000010101)) color_data = 12'b100101110011;
		if(({row_reg, col_reg}==12'b011000010110)) color_data = 12'b100001010010;
		if(({row_reg, col_reg}==12'b011000010111)) color_data = 12'b100001100010;
		if(({row_reg, col_reg}==12'b011000011000)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}>=12'b011000011001) && ({row_reg, col_reg}<12'b011000011100)) color_data = 12'b101001110100;
		if(({row_reg, col_reg}==12'b011000011100)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b011000011101)) color_data = 12'b101101110101;
		if(({row_reg, col_reg}==12'b011000011110)) color_data = 12'b101000100001;
		if(({row_reg, col_reg}==12'b011000011111)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b011000100000) && ({row_reg, col_reg}<12'b011001001100)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b011001001100) && ({row_reg, col_reg}<12'b011001001110)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b011001001110)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=12'b011001001111) && ({row_reg, col_reg}<12'b011001010001)) color_data = 12'b100000010000;
		if(({row_reg, col_reg}==12'b011001010001)) color_data = 12'b011000010000;
		if(({row_reg, col_reg}==12'b011001010010)) color_data = 12'b100001100011;
		if(({row_reg, col_reg}==12'b011001010011)) color_data = 12'b101010010101;
		if(({row_reg, col_reg}==12'b011001010100)) color_data = 12'b100110000100;
		if(({row_reg, col_reg}==12'b011001010101)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==12'b011001010110)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==12'b011001010111)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==12'b011001011000)) color_data = 12'b100001100011;
		if(({row_reg, col_reg}>=12'b011001011001) && ({row_reg, col_reg}<12'b011001011100)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==12'b011001011100)) color_data = 12'b100101110101;
		if(({row_reg, col_reg}==12'b011001011101)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==12'b011001011110)) color_data = 12'b011100010000;
		if(({row_reg, col_reg}==12'b011001011111)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b011001100000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b011001100001) && ({row_reg, col_reg}<12'b011001100101)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b011001100101)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b011001100110) && ({row_reg, col_reg}<12'b011010001101)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b011010001101) && ({row_reg, col_reg}<12'b011010010000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b011010010000)) color_data = 12'b101000010000;
		if(({row_reg, col_reg}==12'b011010010001)) color_data = 12'b011100010000;
		if(({row_reg, col_reg}==12'b011010010010)) color_data = 12'b011000110001;
		if(({row_reg, col_reg}==12'b011010010011)) color_data = 12'b011101100100;
		if(({row_reg, col_reg}==12'b011010010100)) color_data = 12'b011101110100;
		if(({row_reg, col_reg}==12'b011010010101)) color_data = 12'b100110000101;
		if(({row_reg, col_reg}==12'b011010010110)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==12'b011010010111)) color_data = 12'b100110000101;
		if(({row_reg, col_reg}>=12'b011010011000) && ({row_reg, col_reg}<12'b011010011011)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==12'b011010011011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==12'b011010011100)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==12'b011010011101)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==12'b011010011110)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==12'b011010011111)) color_data = 12'b100000110010;
		if(({row_reg, col_reg}==12'b011010100000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}>=12'b011010100001) && ({row_reg, col_reg}<12'b011010100101)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b011010100101)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b011010100110) && ({row_reg, col_reg}<12'b011011010000)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b011011010000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b011011010001)) color_data = 12'b100000100001;
		if(({row_reg, col_reg}==12'b011011010010)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==12'b011011010011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011011010100)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==12'b011011010101)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==12'b011011010110)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}==12'b011011010111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==12'b011011011000)) color_data = 12'b011001100100;
		if(({row_reg, col_reg}>=12'b011011011001) && ({row_reg, col_reg}<12'b011011011011)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==12'b011011011011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011011011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011011011101)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b011011011110)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==12'b011011011111)) color_data = 12'b101010000111;
		if(({row_reg, col_reg}==12'b011011100000)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b011011100001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b011011100010) && ({row_reg, col_reg}<12'b011011100100)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b011011100100) && ({row_reg, col_reg}<12'b011011100110)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b011011100110) && ({row_reg, col_reg}<12'b011100000000)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b011100000000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b011100000001) && ({row_reg, col_reg}<12'b011100001101)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b011100001101)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b011100001110)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b011100001111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b011100010000)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b011100010001)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==12'b011100010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011100010011)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011100010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011100010101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b011100010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011100010111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=12'b011100011000) && ({row_reg, col_reg}<12'b011100011010)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b011100011010)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011100011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011100011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011100011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011100011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011100011111)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==12'b011100100000)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==12'b011100100001)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==12'b011100100010)) color_data = 12'b101100000001;
		if(({row_reg, col_reg}==12'b011100100011)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b011100100100)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b011100100101) && ({row_reg, col_reg}<12'b011101001111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b011101001111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b011101010000)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b011101010001)) color_data = 12'b101001110111;
		if(({row_reg, col_reg}==12'b011101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011101010011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==12'b011101010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011101010101)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}>=12'b011101010110) && ({row_reg, col_reg}<12'b011101011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011101011010)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b011101011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011101011100)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==12'b011101011101)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==12'b011101011110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b011101011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011101100000)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==12'b011101100001)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b011101100010)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b011101100011) && ({row_reg, col_reg}<12'b011110001111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b011110001111)) color_data = 12'b101000000001;
		if(({row_reg, col_reg}==12'b011110010000)) color_data = 12'b100000100010;
		if(({row_reg, col_reg}==12'b011110010001)) color_data = 12'b101001110111;
		if(({row_reg, col_reg}==12'b011110010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011110010011)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b011110010100)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b011110010101)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011110010110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b011110010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011110011000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=12'b011110011001) && ({row_reg, col_reg}<12'b011110011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011110011100)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==12'b011110011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011110011110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b011110011111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b011110100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==12'b011110100001)) color_data = 12'b100000100010;
		if(({row_reg, col_reg}==12'b011110100010)) color_data = 12'b100100000001;

		if(({row_reg, col_reg}>=12'b011110100011) && ({row_reg, col_reg}<12'b011111001111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b011111001111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b011111010000)) color_data = 12'b100100110011;
		if(({row_reg, col_reg}==12'b011111010001)) color_data = 12'b100101100110;
		if(({row_reg, col_reg}==12'b011111010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011111010011)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b011111010100)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==12'b011111010101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=12'b011111010110) && ({row_reg, col_reg}<12'b011111011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011111011010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b011111011011)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b011111011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011111011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011111011110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==12'b011111011111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b011111100000)) color_data = 12'b110010101001;
		if(({row_reg, col_reg}==12'b011111100001)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==12'b011111100010)) color_data = 12'b101000000001;

		if(({row_reg, col_reg}>=12'b011111100011) && ({row_reg, col_reg}<12'b100000001111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b100000001111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b100000010000)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b100000010001)) color_data = 12'b101101110111;
		if(({row_reg, col_reg}==12'b100000010010)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==12'b100000010011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=12'b100000010100) && ({row_reg, col_reg}<12'b100000010110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=12'b100000010110) && ({row_reg, col_reg}<12'b100000011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100000011011)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b100000011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100000011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100000011110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b100000011111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b100000100000)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}==12'b100000100001)) color_data = 12'b100000100010;
		if(({row_reg, col_reg}==12'b100000100010)) color_data = 12'b101000000001;
		if(({row_reg, col_reg}==12'b100000100011)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b100000100100)) color_data = 12'b110000000000;

		if(({row_reg, col_reg}>=12'b100000100101) && ({row_reg, col_reg}<12'b100001001111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b100001001111)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b100001010000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b100001010001)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==12'b100001010010)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==12'b100001010011)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==12'b100001010100)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==12'b100001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100001010110)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=12'b100001010111) && ({row_reg, col_reg}<12'b100001011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100001011001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==12'b100001011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100001011011)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b100001011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001011101)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==12'b100001011110)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b100001011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b100001100000)) color_data = 12'b101001100101;
		if(({row_reg, col_reg}==12'b100001100001)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b100001100010)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b100001100011) && ({row_reg, col_reg}<12'b100010010000)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b100010010000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b100010010001)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b100010010010)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==12'b100010010011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=12'b100010010100) && ({row_reg, col_reg}<12'b100010010110)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==12'b100010010110)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==12'b100010010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}>=12'b100010011000) && ({row_reg, col_reg}<12'b100010011011)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==12'b100010011011)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100010011100)) color_data = 12'b010001010101;
		if(({row_reg, col_reg}==12'b100010011101)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==12'b100010011110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b100010011111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b100010100000)) color_data = 12'b100000110011;
		if(({row_reg, col_reg}==12'b100010100001)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==12'b100010100010)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b100010100011) && ({row_reg, col_reg}<12'b100011010000)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b100011010000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b100011010001)) color_data = 12'b100100010001;
		if(({row_reg, col_reg}==12'b100011010010)) color_data = 12'b011000110011;
		if(({row_reg, col_reg}==12'b100011010011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b100011010100)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==12'b100011010101)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==12'b100011010110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100011010111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100011011000)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==12'b100011011001)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==12'b100011011010)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==12'b100011011011)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==12'b100011011100)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==12'b100011011101)) color_data = 12'b010001100110;
		if(({row_reg, col_reg}==12'b100011011110)) color_data = 12'b010001100101;
		if(({row_reg, col_reg}==12'b100011011111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==12'b100011100000)) color_data = 12'b011100010001;
		if(({row_reg, col_reg}==12'b100011100001)) color_data = 12'b100100000000;

		if(({row_reg, col_reg}>=12'b100011100010) && ({row_reg, col_reg}<12'b100100010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b100100010001)) color_data = 12'b100100010000;
		if(({row_reg, col_reg}==12'b100100010010)) color_data = 12'b011000010001;
		if(({row_reg, col_reg}==12'b100100010011)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==12'b100100010100)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==12'b100100010101)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==12'b100100010110)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==12'b100100010111)) color_data = 12'b001101000100;
		if(({row_reg, col_reg}==12'b100100011000)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==12'b100100011001)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==12'b100100011010)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}==12'b100100011011)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b100100011100)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==12'b100100011101)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==12'b100100011110)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}==12'b100100011111)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==12'b100100100000)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b100100100001)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b100100100010) && ({row_reg, col_reg}<12'b100101010000)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b100101010000) && ({row_reg, col_reg}<12'b100101010010)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b100101010010)) color_data = 12'b011000010000;
		if(({row_reg, col_reg}==12'b100101010011)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==12'b100101010100)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==12'b100101010101)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b100101010110)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==12'b100101010111)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==12'b100101011000)) color_data = 12'b010001100110;
		if(({row_reg, col_reg}==12'b100101011001)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}==12'b100101011010)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}==12'b100101011011)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==12'b100101011100)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==12'b100101011101)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==12'b100101011110)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b100101011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b100101100000)) color_data = 12'b100100010001;

		if(({row_reg, col_reg}>=12'b100101100001) && ({row_reg, col_reg}<12'b100110010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b100110010001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b100110010010)) color_data = 12'b100000010000;
		if(({row_reg, col_reg}==12'b100110010011)) color_data = 12'b100101100101;
		if(({row_reg, col_reg}==12'b100110010100)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}>=12'b100110010101) && ({row_reg, col_reg}<12'b100110010111)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==12'b100110010111)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b100110011000)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==12'b100110011001)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}>=12'b100110011010) && ({row_reg, col_reg}<12'b100110011100)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==12'b100110011100)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b100110011101)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==12'b100110011110)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b100110011111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b100110100000)) color_data = 12'b100100010001;
		if(({row_reg, col_reg}>=12'b100110100001) && ({row_reg, col_reg}<12'b100110100100)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b100110100100)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b100110100101) && ({row_reg, col_reg}<12'b100111010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b100111010001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b100111010010)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==12'b100111010011)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==12'b100111010100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b100111010101)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==12'b100111010110)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==12'b100111010111)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b100111011000)) color_data = 12'b010110001000;
		if(({row_reg, col_reg}==12'b100111011001)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b100111011010)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}>=12'b100111011011) && ({row_reg, col_reg}<12'b100111011101)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==12'b100111011101)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==12'b100111011110)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b100111011111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b100111100000)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b100111100001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b100111100010) && ({row_reg, col_reg}<12'b100111100100)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b100111100100)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b100111100101) && ({row_reg, col_reg}<12'b101000010010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b101000010010)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b101000010011)) color_data = 12'b011100100001;
		if(({row_reg, col_reg}==12'b101000010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b101000010101)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}==12'b101000010110)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}==12'b101000010111)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==12'b101000011000)) color_data = 12'b010110001000;
		if(({row_reg, col_reg}>=12'b101000011001) && ({row_reg, col_reg}<12'b101000011011)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==12'b101000011011)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==12'b101000011100)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}>=12'b101000011101) && ({row_reg, col_reg}<12'b101000011111)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b101000011111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==12'b101000100000)) color_data = 12'b100000010000;
		if(({row_reg, col_reg}==12'b101000100001)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b101000100010) && ({row_reg, col_reg}<12'b101001010010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b101001010010)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b101001010011)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b101001010100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b101001010101)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==12'b101001010110)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==12'b101001010111)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==12'b101001011000)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==12'b101001011001)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==12'b101001011010)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}>=12'b101001011011) && ({row_reg, col_reg}<12'b101001011101)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==12'b101001011101)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==12'b101001011110)) color_data = 12'b100111001010;
		if(({row_reg, col_reg}==12'b101001011111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==12'b101001100000)) color_data = 12'b011100010000;
		if(({row_reg, col_reg}==12'b101001100001)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b101001100010) && ({row_reg, col_reg}<12'b101010010010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b101010010010)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b101010010011)) color_data = 12'b100100100010;
		if(({row_reg, col_reg}==12'b101010010100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=12'b101010010101) && ({row_reg, col_reg}<12'b101010011001)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==12'b101010011001)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==12'b101010011010)) color_data = 12'b010110000111;
		if(({row_reg, col_reg}==12'b101010011011)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}>=12'b101010011100) && ({row_reg, col_reg}<12'b101010011110)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==12'b101010011110)) color_data = 12'b011010011000;
		if(({row_reg, col_reg}==12'b101010011111)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}==12'b101010100000)) color_data = 12'b100000100001;
		if(({row_reg, col_reg}>=12'b101010100001) && ({row_reg, col_reg}<12'b101010100011)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b101010100011) && ({row_reg, col_reg}<12'b101011010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b101011010001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b101011010010)) color_data = 12'b101000000001;
		if(({row_reg, col_reg}==12'b101011010011)) color_data = 12'b011100010001;
		if(({row_reg, col_reg}==12'b101011010100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==12'b101011010101)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}>=12'b101011010110) && ({row_reg, col_reg}<12'b101011011000)) color_data = 12'b101111011100;
		if(({row_reg, col_reg}==12'b101011011000)) color_data = 12'b110011011101;
		if(({row_reg, col_reg}==12'b101011011001)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==12'b101011011010)) color_data = 12'b101111001100;
		if(({row_reg, col_reg}==12'b101011011011)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==12'b101011011100)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b101011011101)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==12'b101011011110)) color_data = 12'b101011001010;
		if(({row_reg, col_reg}==12'b101011011111)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==12'b101011100000)) color_data = 12'b100100110010;
		if(({row_reg, col_reg}==12'b101011100001)) color_data = 12'b101000010000;

		if(({row_reg, col_reg}>=12'b101011100010) && ({row_reg, col_reg}<12'b101100010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b101100010001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b101100010010)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==12'b101100010011)) color_data = 12'b011100110010;
		if(({row_reg, col_reg}==12'b101100010100)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==12'b101100010101)) color_data = 12'b010001010100;
		if(({row_reg, col_reg}==12'b101100010110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==12'b101100010111)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=12'b101100011000) && ({row_reg, col_reg}<12'b101100011010)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b101100011010)) color_data = 12'b101010111001;
		if(({row_reg, col_reg}>=12'b101100011011) && ({row_reg, col_reg}<12'b101100011101)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b101100011101)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b101100011110)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b101100011111)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==12'b101100100000)) color_data = 12'b100000100001;
		if(({row_reg, col_reg}>=12'b101100100001) && ({row_reg, col_reg}<12'b101100100011)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b101100100011) && ({row_reg, col_reg}<12'b101101010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b101101010001)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b101101010010)) color_data = 12'b101101100101;
		if(({row_reg, col_reg}==12'b101101010011)) color_data = 12'b111011001011;
		if(({row_reg, col_reg}==12'b101101010100)) color_data = 12'b110111001011;
		if(({row_reg, col_reg}==12'b101101010101)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==12'b101101010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==12'b101101010111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==12'b101101011000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==12'b101101011001)) color_data = 12'b010101010100;
		if(({row_reg, col_reg}>=12'b101101011010) && ({row_reg, col_reg}<12'b101101011100)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==12'b101101011100)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}>=12'b101101011101) && ({row_reg, col_reg}<12'b101101011111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==12'b101101011111)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==12'b101101100000)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b101101100001)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b101101100010) && ({row_reg, col_reg}<12'b101110010000)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b101110010000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b101110010001)) color_data = 12'b100100010000;
		if(({row_reg, col_reg}==12'b101110010010)) color_data = 12'b111010111010;
		if(({row_reg, col_reg}==12'b101110010011)) color_data = 12'b110111011011;
		if(({row_reg, col_reg}==12'b101110010100)) color_data = 12'b110011011011;
		if(({row_reg, col_reg}==12'b101110010101)) color_data = 12'b111011101100;
		if(({row_reg, col_reg}==12'b101110010110)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==12'b101110010111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==12'b101110011000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==12'b101110011001)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==12'b101110011010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==12'b101110011011)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==12'b101110011100)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==12'b101110011101)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==12'b101110011110)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==12'b101110011111)) color_data = 12'b101001010101;
		if(({row_reg, col_reg}==12'b101110100000)) color_data = 12'b100100010001;

		if(({row_reg, col_reg}>=12'b101110100001) && ({row_reg, col_reg}<12'b101111010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b101111010001)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==12'b101111010010)) color_data = 12'b101001110110;
		if(({row_reg, col_reg}==12'b101111010011)) color_data = 12'b111011001011;
		if(({row_reg, col_reg}==12'b101111010100)) color_data = 12'b110111001010;
		if(({row_reg, col_reg}==12'b101111010101)) color_data = 12'b111011011011;
		if(({row_reg, col_reg}==12'b101111010110)) color_data = 12'b110010001000;
		if(({row_reg, col_reg}==12'b101111010111)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==12'b101111011000)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==12'b101111011001)) color_data = 12'b111010111010;
		if(({row_reg, col_reg}==12'b101111011010)) color_data = 12'b111011011011;
		if(({row_reg, col_reg}==12'b101111011011)) color_data = 12'b110111001010;
		if(({row_reg, col_reg}==12'b101111011100)) color_data = 12'b110110111010;
		if(({row_reg, col_reg}==12'b101111011101)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==12'b101111011110)) color_data = 12'b100001000100;
		if(({row_reg, col_reg}==12'b101111011111)) color_data = 12'b100000100010;
		if(({row_reg, col_reg}==12'b101111100000)) color_data = 12'b100100000000;

		if(({row_reg, col_reg}>=12'b101111100001) && ({row_reg, col_reg}<12'b110000010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b110000010001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b110000010010)) color_data = 12'b011100000000;
		if(({row_reg, col_reg}==12'b110000010011)) color_data = 12'b011100100001;
		if(({row_reg, col_reg}==12'b110000010100)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==12'b110000010101)) color_data = 12'b100101000011;
		if(({row_reg, col_reg}==12'b110000010110)) color_data = 12'b100100110011;
		if(({row_reg, col_reg}==12'b110000010111)) color_data = 12'b100000100010;
		if(({row_reg, col_reg}==12'b110000011000)) color_data = 12'b011100100001;
		if(({row_reg, col_reg}==12'b110000011001)) color_data = 12'b111010111010;
		if(({row_reg, col_reg}==12'b110000011010)) color_data = 12'b110111001011;
		if(({row_reg, col_reg}==12'b110000011011)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==12'b110000011100)) color_data = 12'b110111011011;
		if(({row_reg, col_reg}==12'b110000011101)) color_data = 12'b101110101000;
		if(({row_reg, col_reg}==12'b110000011110)) color_data = 12'b100101100101;
		if(({row_reg, col_reg}==12'b110000011111)) color_data = 12'b011100100001;
		if(({row_reg, col_reg}==12'b110000100000)) color_data = 12'b100100000000;

		if(({row_reg, col_reg}>=12'b110000100001) && ({row_reg, col_reg}<12'b110001010001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b110001010001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b110001010010)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b110001010011)) color_data = 12'b100100010000;
		if(({row_reg, col_reg}==12'b110001010100)) color_data = 12'b100000010000;
		if(({row_reg, col_reg}==12'b110001010101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==12'b110001010110)) color_data = 12'b100100010000;
		if(({row_reg, col_reg}>=12'b110001010111) && ({row_reg, col_reg}<12'b110001011001)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b110001011001)) color_data = 12'b100000110010;
		if(({row_reg, col_reg}==12'b110001011010)) color_data = 12'b101101110110;
		if(({row_reg, col_reg}==12'b110001011011)) color_data = 12'b101110000111;
		if(({row_reg, col_reg}==12'b110001011100)) color_data = 12'b101110010111;
		if(({row_reg, col_reg}==12'b110001011101)) color_data = 12'b110010011000;
		if(({row_reg, col_reg}==12'b110001011110)) color_data = 12'b101001010100;
		if(({row_reg, col_reg}==12'b110001011111)) color_data = 12'b100000010001;
		if(({row_reg, col_reg}==12'b110001100000)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b110001100001) && ({row_reg, col_reg}<12'b110010010010)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b110010010010) && ({row_reg, col_reg}<12'b110010011000)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b110010011000)) color_data = 12'b100100000000;
		if(({row_reg, col_reg}==12'b110010011001)) color_data = 12'b100100010000;
		if(({row_reg, col_reg}>=12'b110010011010) && ({row_reg, col_reg}<12'b110010011100)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}==12'b110010011100)) color_data = 12'b100000010000;
		if(({row_reg, col_reg}==12'b110010011101)) color_data = 12'b100000000000;
		if(({row_reg, col_reg}>=12'b110010011110) && ({row_reg, col_reg}<12'b110010100000)) color_data = 12'b100100000000;

		if(({row_reg, col_reg}>=12'b110010100000) && ({row_reg, col_reg}<12'b110011010111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}>=12'b110011010111) && ({row_reg, col_reg}<12'b110011011100)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}==12'b110011011100)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b110011011101)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b110011011110) && ({row_reg, col_reg}<12'b110100011001)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b110100011001)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b110100011010) && ({row_reg, col_reg}<12'b110100011100)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b110100011100)) color_data = 12'b101000000000;
		if(({row_reg, col_reg}>=12'b110100011101) && ({row_reg, col_reg}<12'b110100011111)) color_data = 12'b101100000000;
		if(({row_reg, col_reg}==12'b110100011111)) color_data = 12'b101000000000;

		if(({row_reg, col_reg}>=12'b110100100000) && ({row_reg, col_reg}<=12'b110100101111)) color_data = 12'b101100000000;
	end
endmodule