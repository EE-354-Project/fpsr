module lebron_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=11'b00000000000) && ({row_reg, col_reg}<11'b00000010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b00000010001)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==11'b00000010010)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==11'b00000010011)) color_data = 12'b111111111110;

		if(({row_reg, col_reg}>=11'b00000010100) && ({row_reg, col_reg}<11'b00001001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b00001001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==11'b00001010000)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}>=11'b00001010001) && ({row_reg, col_reg}<11'b00001010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==11'b00001010011)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==11'b00001010100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==11'b00001010101)) color_data = 12'b111111111110;

		if(({row_reg, col_reg}>=11'b00001010110) && ({row_reg, col_reg}<11'b00010001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b00010001110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==11'b00010001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==11'b00010010000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==11'b00010010001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b00010010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==11'b00010010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==11'b00010010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==11'b00010010101)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==11'b00010010110)) color_data = 12'b111111111110;

		if(({row_reg, col_reg}>=11'b00010010111) && ({row_reg, col_reg}<11'b00011001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b00011001101)) color_data = 12'b110011001011;
		if(({row_reg, col_reg}==11'b00011001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==11'b00011001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00011010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00011010001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==11'b00011010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=11'b00011010011) && ({row_reg, col_reg}<11'b00011010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00011010101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==11'b00011010110)) color_data = 12'b011001010100;

		if(({row_reg, col_reg}>=11'b00011010111) && ({row_reg, col_reg}<11'b00100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b00100001101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==11'b00100001110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==11'b00100001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b00100010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b00100010001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00100010010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=11'b00100010011) && ({row_reg, col_reg}<11'b00100010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00100010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00100010110)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==11'b00100010111)) color_data = 12'b110010111011;

		if(({row_reg, col_reg}>=11'b00100011000) && ({row_reg, col_reg}<11'b00101001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b00101001101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b00101001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b00101001111)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==11'b00101010000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00101010001)) color_data = 12'b011000110010;
		if(({row_reg, col_reg}==11'b00101010010)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=11'b00101010011) && ({row_reg, col_reg}<11'b00101010101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b00101010101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00101010110)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==11'b00101010111)) color_data = 12'b101010011000;

		if(({row_reg, col_reg}>=11'b00101011000) && ({row_reg, col_reg}<11'b00110001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b00110001101)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==11'b00110001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==11'b00110001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00110010001)) color_data = 12'b011000110010;
		if(({row_reg, col_reg}==11'b00110010010)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b00110010011)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b00110010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00110010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b00110010110)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==11'b00110010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==11'b00110011000)) color_data = 12'b111111111110;

		if(({row_reg, col_reg}>=11'b00110011001) && ({row_reg, col_reg}<11'b00111001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b00111001100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==11'b00111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=11'b00111001110) && ({row_reg, col_reg}<11'b00111010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00111010000)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==11'b00111010001)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==11'b00111010010)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==11'b00111010011)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}>=11'b00111010100) && ({row_reg, col_reg}<11'b00111010110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b00111010110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b00111010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b00111011000)) color_data = 12'b110010111011;

		if(({row_reg, col_reg}>=11'b00111011001) && ({row_reg, col_reg}<11'b01000001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b01000001100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b01000001101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==11'b01000001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=11'b01000001111) && ({row_reg, col_reg}<11'b01000010001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01000010001)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==11'b01000010010)) color_data = 12'b011000110010;
		if(({row_reg, col_reg}==11'b01000010011)) color_data = 12'b010000100000;
		if(({row_reg, col_reg}==11'b01000010100)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==11'b01000010101)) color_data = 12'b010101000010;
		if(({row_reg, col_reg}==11'b01000010110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01000010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==11'b01000011000)) color_data = 12'b101010011000;

		if(({row_reg, col_reg}>=11'b01000011001) && ({row_reg, col_reg}<11'b01001001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b01001001100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b01001001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b01001001110)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01001001111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01001010000)) color_data = 12'b011000110010;
		if(({row_reg, col_reg}==11'b01001010001)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==11'b01001010010)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b01001010011)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==11'b01001010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01001010101)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01001010110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01001010111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b01001011000)) color_data = 12'b100110001000;

		if(({row_reg, col_reg}>=11'b01001011001) && ({row_reg, col_reg}<11'b01010001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b01010001100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==11'b01010001101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==11'b01010001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01010001111)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01010010000)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==11'b01010010001)) color_data = 12'b011000110010;
		if(({row_reg, col_reg}==11'b01010010010)) color_data = 12'b010100100001;
		if(({row_reg, col_reg}==11'b01010010011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01010010100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01010010101)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b01010010110)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b01010010111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==11'b01010011000)) color_data = 12'b101110101010;

		if(({row_reg, col_reg}>=11'b01010011001) && ({row_reg, col_reg}<11'b01011001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b01011001100)) color_data = 12'b111111101110;
		if(({row_reg, col_reg}==11'b01011001101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==11'b01011001110)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==11'b01011001111)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01011010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01011010001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b01011010010)) color_data = 12'b011000110010;
		if(({row_reg, col_reg}==11'b01011010011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b01011010100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b01011010101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b01011010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01011010111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==11'b01011011000)) color_data = 12'b111011011101;

		if(({row_reg, col_reg}>=11'b01011011001) && ({row_reg, col_reg}<11'b01100001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b01100001101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==11'b01100001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==11'b01100001111)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==11'b01100010000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01100010001)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==11'b01100010010)) color_data = 12'b101110011000;
		if(({row_reg, col_reg}==11'b01100010011)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}>=11'b01100010100) && ({row_reg, col_reg}<11'b01100010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01100010110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==11'b01100010111)) color_data = 12'b001100100010;

		if(({row_reg, col_reg}>=11'b01100011000) && ({row_reg, col_reg}<11'b01101001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b01101001101)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==11'b01101001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==11'b01101001111)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}>=11'b01101010000) && ({row_reg, col_reg}<11'b01101010010)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==11'b01101010010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101010011)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b01101010100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b01101010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==11'b01101010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==11'b01101010111)) color_data = 12'b001100110011;

		if(({row_reg, col_reg}>=11'b01101011000) && ({row_reg, col_reg}<11'b01110001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b01110001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=11'b01110001110) && ({row_reg, col_reg}<11'b01110010000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==11'b01110010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==11'b01110010001)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==11'b01110010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==11'b01110010011)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==11'b01110010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==11'b01110010101)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==11'b01110010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==11'b01110010111)) color_data = 12'b011101100110;

		if(({row_reg, col_reg}>=11'b01110011000) && ({row_reg, col_reg}<11'b01111001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b01111001101)) color_data = 12'b110111001100;
		if(({row_reg, col_reg}>=11'b01111001110) && ({row_reg, col_reg}<11'b01111010001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==11'b01111010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}==11'b01111010010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==11'b01111010011)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=11'b01111010100) && ({row_reg, col_reg}<11'b01111010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==11'b01111010111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=11'b01111011000) && ({row_reg, col_reg}<11'b10000001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b10000001110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=11'b10000001111) && ({row_reg, col_reg}<11'b10000010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==11'b10000010110)) color_data = 12'b010001000100;

		if(({row_reg, col_reg}>=11'b10000010111) && ({row_reg, col_reg}<11'b10001001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=11'b10001001010) && ({row_reg, col_reg}<11'b10001001101)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==11'b10001001101)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==11'b10001001110)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b10001001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b10001010000)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==11'b10001010001)) color_data = 12'b000100010000;
		if(({row_reg, col_reg}>=11'b10001010010) && ({row_reg, col_reg}<11'b10001010100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==11'b10001010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==11'b10001010101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==11'b10001010110)) color_data = 12'b001100110010;
		if(({row_reg, col_reg}==11'b10001010111)) color_data = 12'b010001000011;
		if(({row_reg, col_reg}==11'b10001011000)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b10001011001)) color_data = 12'b111111101101;

		if(({row_reg, col_reg}>=11'b10001011010) && ({row_reg, col_reg}<11'b10010001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b10010001010)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==11'b10010001011)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}>=11'b10010001100) && ({row_reg, col_reg}<11'b10010001110)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==11'b10010001110)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b10010001111)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b10010010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}>=11'b10010010001) && ({row_reg, col_reg}<11'b10010010100)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b10010010100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==11'b10010010101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b10010010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b10010010111)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==11'b10010011000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==11'b10010011001)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==11'b10010011010)) color_data = 12'b110110111001;
		if(({row_reg, col_reg}==11'b10010011011)) color_data = 12'b111111101011;
		if(({row_reg, col_reg}==11'b10010011100)) color_data = 12'b111111111110;

		if(({row_reg, col_reg}>=11'b10010011101) && ({row_reg, col_reg}<11'b10011000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=11'b10011000111) && ({row_reg, col_reg}<11'b10011001001)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==11'b10011001001)) color_data = 12'b111011011011;
		if(({row_reg, col_reg}==11'b10011001010)) color_data = 12'b110010100111;
		if(({row_reg, col_reg}==11'b10011001011)) color_data = 12'b100101110100;
		if(({row_reg, col_reg}==11'b10011001100)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==11'b10011001101)) color_data = 12'b010101000001;
		if(({row_reg, col_reg}==11'b10011001110)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==11'b10011001111)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==11'b10011010000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==11'b10011010001)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==11'b10011010010)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==11'b10011010011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b10011010100)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b10011010101)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=11'b10011010110) && ({row_reg, col_reg}<11'b10011011001)) color_data = 12'b010100110001;
		if(({row_reg, col_reg}==11'b10011011001)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==11'b10011011010)) color_data = 12'b100101110011;
		if(({row_reg, col_reg}==11'b10011011011)) color_data = 12'b100001110011;
		if(({row_reg, col_reg}==11'b10011011100)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==11'b10011011101)) color_data = 12'b111111111110;

		if(({row_reg, col_reg}>=11'b10011011110) && ({row_reg, col_reg}<11'b10100000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b10100000111)) color_data = 12'b111111011101;
		if(({row_reg, col_reg}==11'b10100001000)) color_data = 12'b110010110111;
		if(({row_reg, col_reg}==11'b10100001001)) color_data = 12'b101110100101;
		if(({row_reg, col_reg}==11'b10100001010)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==11'b10100001011)) color_data = 12'b110110110101;
		if(({row_reg, col_reg}==11'b10100001100)) color_data = 12'b100101110011;
		if(({row_reg, col_reg}>=11'b10100001101) && ({row_reg, col_reg}<11'b10100001111)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==11'b10100001111)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==11'b10100010000)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==11'b10100010001)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}>=11'b10100010010) && ({row_reg, col_reg}<11'b10100010100)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=11'b10100010100) && ({row_reg, col_reg}<11'b10100010110)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}>=11'b10100010110) && ({row_reg, col_reg}<11'b10100011000)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==11'b10100011000)) color_data = 12'b101110010100;
		if(({row_reg, col_reg}==11'b10100011001)) color_data = 12'b110110110111;
		if(({row_reg, col_reg}==11'b10100011010)) color_data = 12'b101010000011;
		if(({row_reg, col_reg}==11'b10100011011)) color_data = 12'b010100110000;
		if(({row_reg, col_reg}==11'b10100011100)) color_data = 12'b001100100000;
		if(({row_reg, col_reg}==11'b10100011101)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b10100011110)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==11'b10100011111)) color_data = 12'b111111011101;

		if(({row_reg, col_reg}>=11'b10100100000) && ({row_reg, col_reg}<11'b10101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b10101000110)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==11'b10101000111)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==11'b10101001000)) color_data = 12'b100101110011;
		if(({row_reg, col_reg}==11'b10101001001)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==11'b10101001010)) color_data = 12'b110110110010;
		if(({row_reg, col_reg}==11'b10101001011)) color_data = 12'b111011000011;
		if(({row_reg, col_reg}==11'b10101001100)) color_data = 12'b110110110101;
		if(({row_reg, col_reg}==11'b10101001101)) color_data = 12'b100101110011;
		if(({row_reg, col_reg}==11'b10101001110)) color_data = 12'b011101000001;
		if(({row_reg, col_reg}==11'b10101001111)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==11'b10101010000)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}>=11'b10101010001) && ({row_reg, col_reg}<11'b10101010011)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==11'b10101010011)) color_data = 12'b100101100011;
		if(({row_reg, col_reg}==11'b10101010100)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}==11'b10101010101)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==11'b10101010110)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==11'b10101010111)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}==11'b10101011000)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==11'b10101011001)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==11'b10101011010)) color_data = 12'b111111000110;
		if(({row_reg, col_reg}==11'b10101011011)) color_data = 12'b110110100110;
		if(({row_reg, col_reg}==11'b10101011100)) color_data = 12'b100001100100;
		if(({row_reg, col_reg}==11'b10101011101)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b10101011110)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==11'b10101011111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b10101100000)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==11'b10101100001)) color_data = 12'b111111111110;

		if(({row_reg, col_reg}>=11'b10101100010) && ({row_reg, col_reg}<11'b10110000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b10110000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==11'b10110000101)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==11'b10110000110)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==11'b10110000111)) color_data = 12'b011101010010;
		if(({row_reg, col_reg}==11'b10110001000)) color_data = 12'b100110000011;
		if(({row_reg, col_reg}==11'b10110001001)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==11'b10110001010)) color_data = 12'b111011000010;
		if(({row_reg, col_reg}==11'b10110001011)) color_data = 12'b111011000001;
		if(({row_reg, col_reg}==11'b10110001100)) color_data = 12'b111011000011;
		if(({row_reg, col_reg}==11'b10110001101)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==11'b10110001110)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}==11'b10110001111)) color_data = 12'b100001010010;
		if(({row_reg, col_reg}==11'b10110010000)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==11'b10110010001)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}>=11'b10110010010) && ({row_reg, col_reg}<11'b10110010100)) color_data = 12'b100001100011;
		if(({row_reg, col_reg}==11'b10110010100)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==11'b10110010101)) color_data = 12'b100001010010;
		if(({row_reg, col_reg}==11'b10110010110)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==11'b10110010111)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==11'b10110011000)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==11'b10110011001)) color_data = 12'b110110100010;
		if(({row_reg, col_reg}==11'b10110011010)) color_data = 12'b111010110100;
		if(({row_reg, col_reg}==11'b10110011011)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==11'b10110011100)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==11'b10110011101)) color_data = 12'b011101100011;
		if(({row_reg, col_reg}>=11'b10110011110) && ({row_reg, col_reg}<11'b10110100000)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b10110100000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==11'b10110100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b10110100010)) color_data = 12'b111111101110;

		if(({row_reg, col_reg}>=11'b10110100011) && ({row_reg, col_reg}<11'b10111000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b10111000010)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==11'b10111000011)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==11'b10111000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b10111000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b10111000110)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==11'b10111000111)) color_data = 12'b100001100010;
		if(({row_reg, col_reg}==11'b10111001000)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==11'b10111001001)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==11'b10111001010)) color_data = 12'b111111010011;
		if(({row_reg, col_reg}==11'b10111001011)) color_data = 12'b111111010001;
		if(({row_reg, col_reg}==11'b10111001100)) color_data = 12'b111111000011;
		if(({row_reg, col_reg}==11'b10111001101)) color_data = 12'b111111010101;
		if(({row_reg, col_reg}==11'b10111001110)) color_data = 12'b111111000110;
		if(({row_reg, col_reg}==11'b10111001111)) color_data = 12'b110110100101;
		if(({row_reg, col_reg}==11'b10111010000)) color_data = 12'b101110000100;
		if(({row_reg, col_reg}==11'b10111010001)) color_data = 12'b100101110010;
		if(({row_reg, col_reg}==11'b10111010010)) color_data = 12'b100001100001;
		if(({row_reg, col_reg}==11'b10111010011)) color_data = 12'b100101110010;
		if(({row_reg, col_reg}==11'b10111010100)) color_data = 12'b101001110011;
		if(({row_reg, col_reg}==11'b10111010101)) color_data = 12'b110010100101;
		if(({row_reg, col_reg}==11'b10111010110)) color_data = 12'b111011000111;
		if(({row_reg, col_reg}==11'b10111010111)) color_data = 12'b110010100011;
		if(({row_reg, col_reg}==11'b10111011000)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==11'b10111011001)) color_data = 12'b110010010001;
		if(({row_reg, col_reg}==11'b10111011010)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==11'b10111011011)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==11'b10111011100)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==11'b10111011101)) color_data = 12'b100001100011;
		if(({row_reg, col_reg}==11'b10111011110)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}>=11'b10111011111) && ({row_reg, col_reg}<11'b10111100001)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b10111100001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==11'b10111100010)) color_data = 12'b011001010101;

		if(({row_reg, col_reg}>=11'b10111100011) && ({row_reg, col_reg}<11'b11000000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b11000000010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==11'b11000000011)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==11'b11000000100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b11000000101)) color_data = 12'b011001000010;
		if(({row_reg, col_reg}==11'b11000000110)) color_data = 12'b011101000010;
		if(({row_reg, col_reg}==11'b11000000111)) color_data = 12'b100001010010;
		if(({row_reg, col_reg}==11'b11000001000)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==11'b11000001001)) color_data = 12'b111011000111;
		if(({row_reg, col_reg}==11'b11000001010)) color_data = 12'b111111010100;
		if(({row_reg, col_reg}==11'b11000001011)) color_data = 12'b111111010011;
		if(({row_reg, col_reg}==11'b11000001100)) color_data = 12'b111111010100;
		if(({row_reg, col_reg}>=11'b11000001101) && ({row_reg, col_reg}<11'b11000001111)) color_data = 12'b111011000011;
		if(({row_reg, col_reg}==11'b11000001111)) color_data = 12'b111111010100;
		if(({row_reg, col_reg}==11'b11000010000)) color_data = 12'b111111010101;
		if(({row_reg, col_reg}==11'b11000010001)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==11'b11000010010)) color_data = 12'b110110110100;
		if(({row_reg, col_reg}==11'b11000010011)) color_data = 12'b110111000100;
		if(({row_reg, col_reg}==11'b11000010100)) color_data = 12'b111011000100;
		if(({row_reg, col_reg}==11'b11000010101)) color_data = 12'b111111010101;
		if(({row_reg, col_reg}==11'b11000010110)) color_data = 12'b111011000100;
		if(({row_reg, col_reg}==11'b11000010111)) color_data = 12'b101010000001;
		if(({row_reg, col_reg}==11'b11000011000)) color_data = 12'b101010000010;
		if(({row_reg, col_reg}==11'b11000011001)) color_data = 12'b101001110010;
		if(({row_reg, col_reg}==11'b11000011010)) color_data = 12'b101001110001;
		if(({row_reg, col_reg}==11'b11000011011)) color_data = 12'b110010100100;
		if(({row_reg, col_reg}==11'b11000011100)) color_data = 12'b101110010110;
		if(({row_reg, col_reg}==11'b11000011101)) color_data = 12'b100101110101;
		if(({row_reg, col_reg}==11'b11000011110)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==11'b11000011111)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==11'b11000100000)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b11000100001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b11000100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b11000100011)) color_data = 12'b101110111010;

		if(({row_reg, col_reg}>=11'b11000100100) && ({row_reg, col_reg}<11'b11001000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b11001000001)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==11'b11001000010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b11001000011)) color_data = 12'b011001010011;
		if(({row_reg, col_reg}==11'b11001000100)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b11001000101)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}>=11'b11001000110) && ({row_reg, col_reg}<11'b11001001000)) color_data = 12'b100001010011;
		if(({row_reg, col_reg}==11'b11001001000)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==11'b11001001001)) color_data = 12'b110111000111;
		if(({row_reg, col_reg}==11'b11001001010)) color_data = 12'b111111010101;
		if(({row_reg, col_reg}==11'b11001001011)) color_data = 12'b110110110010;
		if(({row_reg, col_reg}==11'b11001001100)) color_data = 12'b110010100001;
		if(({row_reg, col_reg}==11'b11001001101)) color_data = 12'b110110110001;
		if(({row_reg, col_reg}>=11'b11001001110) && ({row_reg, col_reg}<11'b11001010000)) color_data = 12'b111111010010;
		if(({row_reg, col_reg}==11'b11001010000)) color_data = 12'b111111010011;
		if(({row_reg, col_reg}==11'b11001010001)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}==11'b11001010010)) color_data = 12'b111011000100;
		if(({row_reg, col_reg}>=11'b11001010011) && ({row_reg, col_reg}<11'b11001010110)) color_data = 12'b111111010011;
		if(({row_reg, col_reg}==11'b11001010110)) color_data = 12'b111011010011;
		if(({row_reg, col_reg}==11'b11001010111)) color_data = 12'b110110110010;
		if(({row_reg, col_reg}==11'b11001011000)) color_data = 12'b101110000010;
		if(({row_reg, col_reg}==11'b11001011001)) color_data = 12'b101110000011;
		if(({row_reg, col_reg}==11'b11001011010)) color_data = 12'b110010010010;
		if(({row_reg, col_reg}==11'b11001011011)) color_data = 12'b111010110101;
		if(({row_reg, col_reg}==11'b11001011100)) color_data = 12'b110110110111;
		if(({row_reg, col_reg}==11'b11001011101)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==11'b11001011110)) color_data = 12'b100001100011;
		if(({row_reg, col_reg}==11'b11001011111)) color_data = 12'b100001100100;
		if(({row_reg, col_reg}==11'b11001100000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b11001100001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==11'b11001100010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==11'b11001100011)) color_data = 12'b011101100101;

		if(({row_reg, col_reg}>=11'b11001100100) && ({row_reg, col_reg}<11'b11010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==11'b11010000001)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==11'b11010000010)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==11'b11010000011)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==11'b11010000100)) color_data = 12'b011101010100;
		if(({row_reg, col_reg}==11'b11010000101)) color_data = 12'b100001010100;
		if(({row_reg, col_reg}==11'b11010000110)) color_data = 12'b100101010011;
		if(({row_reg, col_reg}==11'b11010000111)) color_data = 12'b100001010010;
		if(({row_reg, col_reg}==11'b11010001000)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}==11'b11010001001)) color_data = 12'b111011001000;
		if(({row_reg, col_reg}==11'b11010001010)) color_data = 12'b110010100100;
		if(({row_reg, col_reg}==11'b11010001011)) color_data = 12'b100001100000;
		if(({row_reg, col_reg}==11'b11010001100)) color_data = 12'b110010100010;
		if(({row_reg, col_reg}==11'b11010001101)) color_data = 12'b111111010011;
		if(({row_reg, col_reg}>=11'b11010001110) && ({row_reg, col_reg}<11'b11010010011)) color_data = 12'b111111010010;
		if(({row_reg, col_reg}>=11'b11010010011) && ({row_reg, col_reg}<11'b11010011000)) color_data = 12'b111111010011;
		if(({row_reg, col_reg}==11'b11010011000)) color_data = 12'b110110110011;
		if(({row_reg, col_reg}>=11'b11010011001) && ({row_reg, col_reg}<11'b11010011011)) color_data = 12'b111010110011;
		if(({row_reg, col_reg}==11'b11010011011)) color_data = 12'b111111010101;
		if(({row_reg, col_reg}==11'b11010011100)) color_data = 12'b111011000111;
		if(({row_reg, col_reg}==11'b11010011101)) color_data = 12'b101010000101;
		if(({row_reg, col_reg}>=11'b11010011110) && ({row_reg, col_reg}<11'b11010100000)) color_data = 12'b100001100011;
		if(({row_reg, col_reg}==11'b11010100000)) color_data = 12'b011101010011;
		if(({row_reg, col_reg}==11'b11010100001)) color_data = 12'b010101000011;
		if(({row_reg, col_reg}==11'b11010100010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==11'b11010100011)) color_data = 12'b001100100010;

		if(({row_reg, col_reg}>=11'b11010100100) && ({row_reg, col_reg}<=11'b11010100100)) color_data = 12'b111111101110;
	end
endmodule